module activation(
    input activation_type,
    input enable_activation,
    input in_data_available,
    input [`MAT_MUL_SIZE*`DWIDTH-1:0] inp_data,
    output [`MAT_MUL_SIZE*`DWIDTH-1:0] out_data,
    output out_data_available,
    input [`MASK_WIDTH-1:0] validity_mask,
    output done_activation,
    input clk,
    input reset
);

reg  finish_activation;
reg  out_data_valid;
reg  [`MAT_MUL_SIZE*`DWIDTH-1:0] out_activation;
integer i;

reg [3:0] address[`MAT_MUL_SIZE-1:0];
reg [7:0] data_slope[`MAT_MUL_SIZE-1:0];
reg [7:0] data_intercept[`MAT_MUL_SIZE-1:0];

// If the activation block is not enabled, just forward the input data
assign out_data             = enable_activation ? out_activation    : inp_data;
assign done_activation      = enable_activation ? finish_activation : 1'b1;
assign out_data_available   = enable_activation ? out_data_valid    : in_data_available;

always @(posedge clk) begin
    if (reset) begin
      out_activation   <= {`MAT_MUL_SIZE*`DWIDTH-1{1'b0}};
      finish_activation<= 1'b0;
      out_data_valid   <= 1'b0;
    end
    else begin
       if(in_data_available) begin
           for (i = 0; i < `MAT_MUL_SIZE; i=i+1) begin
               if(activation_type==1'b1) begin // tanH
                    out_activation[i*`DWIDTH +:`DWIDTH] <= data_slope[i] * inp_data[i*`DWIDTH +:`DWIDTH] + data_intercept[i];
               end
               else begin // ReLU
                    out_activation[i*`DWIDTH +:`DWIDTH] <= inp_data[i*`DWIDTH-1] ? {`DWIDTH{1'b0}} : inp_data[i*`DWIDTH +:`DWIDTH];
               end
           end 
           finish_activation<= 1'b1;
           out_data_valid   <= 1'b1;
       end
       else begin
           out_activation   <= {`MAT_MUL_SIZE*`DWIDTH-1{1'b0}};
           finish_activation<= 1'b0;
           out_data_valid   <= 1'b0;
       end
    end
end

//Our equation of tanh is Y=AX+B
//A is the slope and B is the intercept.
//We store A in one LUT and B in another.
//LUT for the slope
always @(address) begin
    for (i = 0; i < `MAT_MUL_SIZE; i=i+1) begin
    case (address[i])
      4'b0000: data_slope[i][7:0] = 8'd0;
      4'b0001: data_slope[i][7:0] = 8'd0;
      4'b0010: data_slope[i][7:0] = 8'd2;
      4'b0011: data_slope[i][7:0] = 8'd3;
      4'b0100: data_slope[i][7:0] = 8'd4;
      4'b0101: data_slope[i][7:0] = 8'd0;
      4'b0110: data_slope[i][7:0] = 8'd4;
      4'b0111: data_slope[i][7:0] = 8'd3;
      4'b1000: data_slope[i][7:0] = 8'd2;
      4'b1001: data_slope[i][7:0] = 8'd0;
      4'b1010: data_slope[i][7:0] = 8'd0;
      default: data_slope[i][7:0] = 8'd0;
    endcase  
    end
end

//LUT for the intercept
always @(address) begin
    for (i = 0; i < `MAT_MUL_SIZE; i=i+1) begin
    case (address[i])
      4'b0000: data_intercept[i][7:0] = 8'd127;
      4'b0001: data_intercept[i][7:0] = 8'd99;
      4'b0010: data_intercept[i][7:0] = 8'd46;
      4'b0011: data_intercept[i][7:0] = 8'd18;
      4'b0100: data_intercept[i][7:0] = 8'd0;
      4'b0101: data_intercept[i][7:0] = 8'd0;
      4'b0110: data_intercept[i][7:0] = 8'd0;
      4'b0111: data_intercept[i][7:0] = -8'd18;
      4'b1000: data_intercept[i][7:0] = -8'd46;
      4'b1001: data_intercept[i][7:0] = -8'd99;
      4'b1010: data_intercept[i][7:0] = -8'd127;
      default: data_intercept[i][7:0] = 8'd0;
    endcase  
    end
end

//Logic to find address
always @(inp_data) begin
    for (i = 0; i < `MAT_MUL_SIZE; i=i+1) begin
        if((inp_data[i*`DWIDTH +:`DWIDTH])>=90) begin
           address[i][3:0] = 4'b0000;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=39 && (inp_data[i*`DWIDTH +:`DWIDTH])<90) begin
           address[i][3:0] = 4'b0001;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=28 && (inp_data[i*`DWIDTH +:`DWIDTH])<39) begin
           address[i][3:0] = 4'b0010;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=16 && (inp_data[i*`DWIDTH +:`DWIDTH])<28) begin
           address[i][3:0] = 4'b0011;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=1 && (inp_data[i*`DWIDTH +:`DWIDTH])<16) begin
           address[i][3:0] = 4'b0100;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])==0) begin
           address[i][3:0] = 4'b0101;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-16 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-1) begin
           address[i][3:0] = 4'b0110;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-28 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-16) begin
           address[i][3:0] = 4'b0111;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-39 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-28) begin
           address[i][3:0] = 4'b1000;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-90 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-39) begin
           address[i][3:0] = 4'b1001;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])<=-90) begin
           address[i][3:0] = 4'b1010;
        end
        else begin
           address[i][3:0] = 4'b0101;
        end
    end
end

//Adding a dummy signal to use validity_mask input, to make ODIN happy
//TODO: Need to correctly use validity_mask
wire [`MASK_WIDTH-1:0] dummy;
assign dummy = validity_mask;

// generate multiple ReLU block based on the MAT_MUL_SIZE
//genvar i;
//generate 
//  for (i = 1; i <= `MAT_MUL_SIZE; i = i + 1) begin : loop_gen_ReLU
//        ReLU ReLUinst (.inp_data(inp_data[i*`DWIDTH-1 -:`DWIDTH]), .out_data(temp[i*`DWIDTH-1 -:`DWIDTH]));
//  end
//endgenerate

endmodule

//module ReLU(
//    input [`DWIDTH-1:0] inp_data,
//    output[`DWIDTH-1:0] out_data
//);
//
//assign out_data = inp_data[`DWIDTH-1] ? {`DWIDTH{1'b0}} : inp_data;
//
//endmodule
