
`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020-07-26 21:33:35.015511
// Design Name: 
// Module Name: matmul_32x32_systolic
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module matmul_32x32_systolic(
 clk,
 reset,
 pe_reset,
 start_mat_mul,
 done_mat_mul,
 address_mat_a,
 address_mat_b,
 address_mat_c,
 address_stride_a,
 address_stride_b,
 address_stride_c,
 a_data,
 b_data,
 a_data_in, //Data values coming in from previous matmul - systolic connections
 b_data_in,
 c_data_in, //Data values coming in from previous matmul - systolic shifting
 c_data_out, //Data values going out to next matmul - systolic shifting
 a_data_out,
 b_data_out,
 a_addr,
 b_addr,
 c_addr,
 c_data_available,

 validity_mask_a_rows,
 validity_mask_a_cols_b_rows,
 validity_mask_b_cols,
  
final_mat_mul_size,
  
 a_loc,
 b_loc
);

 input clk;
 input reset;
 input pe_reset;
 input start_mat_mul;
 output done_mat_mul;
 input [`AWIDTH-1:0] address_mat_a;
 input [`AWIDTH-1:0] address_mat_b;
 input [`AWIDTH-1:0] address_mat_c;
 input [`ADDR_STRIDE_WIDTH-1:0] address_stride_a;
 input [`ADDR_STRIDE_WIDTH-1:0] address_stride_b;
 input [`ADDR_STRIDE_WIDTH-1:0] address_stride_c;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_in;
 output [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out;
 output [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data_out;
 output [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data_out;
 output [`AWIDTH-1:0] a_addr;
 output [`AWIDTH-1:0] b_addr;
 output [`AWIDTH-1:0] c_addr;
 output c_data_available;

 input [`MASK_WIDTH-1:0] validity_mask_a_rows;
 input [`MASK_WIDTH-1:0] validity_mask_a_cols_b_rows;
 input [`MASK_WIDTH-1:0] validity_mask_b_cols;

//7:0 is okay here. We aren't going to make a matmul larger than 128x128
//In fact, these will get optimized out by the synthesis tool, because
//we hardcode them at the instantiation level.
 input [7:0] final_mat_mul_size;
  
 input [7:0] a_loc;
 input [7:0] b_loc;

//////////////////////////////////////////////////////////////////////////
// Logic for clock counting and when to assert done
//////////////////////////////////////////////////////////////////////////

reg done_mat_mul;
//This is 7 bits because the expectation is that clock count will be pretty
//small. For large matmuls, this will need to increased to have more bits.
//In general, a systolic multiplier takes 4*N-2+P cycles, where N is the size 
//of the matmul and P is the number of pipleine stages in the MAC block.
reg [7:0] clk_cnt;

//Finding out number of cycles to assert matmul done.
//When we have to save the outputs to accumulators, then we don't need to
//shift out data. So, we can assert done_mat_mul early.
//In the normal case, we have to include the time to shift out the results. 
//Note: the count expression used to contain "4*final_mat_mul_size", but 
//to avoid multiplication, we now use "final_mat_mul_size<<2"
wire [7:0] clk_cnt_for_done;

assign clk_cnt_for_done = 
                          ((final_mat_mul_size<<2) - 2 + `NUM_CYCLES_IN_MAC);  
    
always @(posedge clk) begin
  if (reset || ~start_mat_mul) begin
    clk_cnt <= 0;
    done_mat_mul <= 0;
  end
  else if (clk_cnt == clk_cnt_for_done) begin
    done_mat_mul <= 1;
    clk_cnt <= clk_cnt + 1;

  end
  else if (done_mat_mul == 0) begin
    clk_cnt <= clk_cnt + 1;

  end    
  else begin
    done_mat_mul <= 0;
    clk_cnt <= clk_cnt + 1;
  end
end
wire [`DWIDTH-1:0] a0_data;
wire [`DWIDTH-1:0] a1_data;
wire [`DWIDTH-1:0] a2_data;
wire [`DWIDTH-1:0] a3_data;
wire [`DWIDTH-1:0] a4_data;
wire [`DWIDTH-1:0] a5_data;
wire [`DWIDTH-1:0] a6_data;
wire [`DWIDTH-1:0] a7_data;
wire [`DWIDTH-1:0] a8_data;
wire [`DWIDTH-1:0] a9_data;
wire [`DWIDTH-1:0] a10_data;
wire [`DWIDTH-1:0] a11_data;
wire [`DWIDTH-1:0] a12_data;
wire [`DWIDTH-1:0] a13_data;
wire [`DWIDTH-1:0] a14_data;
wire [`DWIDTH-1:0] a15_data;
wire [`DWIDTH-1:0] a16_data;
wire [`DWIDTH-1:0] a17_data;
wire [`DWIDTH-1:0] a18_data;
wire [`DWIDTH-1:0] a19_data;
wire [`DWIDTH-1:0] a20_data;
wire [`DWIDTH-1:0] a21_data;
wire [`DWIDTH-1:0] a22_data;
wire [`DWIDTH-1:0] a23_data;
wire [`DWIDTH-1:0] a24_data;
wire [`DWIDTH-1:0] a25_data;
wire [`DWIDTH-1:0] a26_data;
wire [`DWIDTH-1:0] a27_data;
wire [`DWIDTH-1:0] a28_data;
wire [`DWIDTH-1:0] a29_data;
wire [`DWIDTH-1:0] a30_data;
wire [`DWIDTH-1:0] a31_data;
wire [`DWIDTH-1:0] b0_data;
wire [`DWIDTH-1:0] b1_data;
wire [`DWIDTH-1:0] b2_data;
wire [`DWIDTH-1:0] b3_data;
wire [`DWIDTH-1:0] b4_data;
wire [`DWIDTH-1:0] b5_data;
wire [`DWIDTH-1:0] b6_data;
wire [`DWIDTH-1:0] b7_data;
wire [`DWIDTH-1:0] b8_data;
wire [`DWIDTH-1:0] b9_data;
wire [`DWIDTH-1:0] b10_data;
wire [`DWIDTH-1:0] b11_data;
wire [`DWIDTH-1:0] b12_data;
wire [`DWIDTH-1:0] b13_data;
wire [`DWIDTH-1:0] b14_data;
wire [`DWIDTH-1:0] b15_data;
wire [`DWIDTH-1:0] b16_data;
wire [`DWIDTH-1:0] b17_data;
wire [`DWIDTH-1:0] b18_data;
wire [`DWIDTH-1:0] b19_data;
wire [`DWIDTH-1:0] b20_data;
wire [`DWIDTH-1:0] b21_data;
wire [`DWIDTH-1:0] b22_data;
wire [`DWIDTH-1:0] b23_data;
wire [`DWIDTH-1:0] b24_data;
wire [`DWIDTH-1:0] b25_data;
wire [`DWIDTH-1:0] b26_data;
wire [`DWIDTH-1:0] b27_data;
wire [`DWIDTH-1:0] b28_data;
wire [`DWIDTH-1:0] b29_data;
wire [`DWIDTH-1:0] b30_data;
wire [`DWIDTH-1:0] b31_data;
wire [`DWIDTH-1:0] a1_data_delayed_1;
wire [`DWIDTH-1:0] a2_data_delayed_1;
wire [`DWIDTH-1:0] a2_data_delayed_2;
wire [`DWIDTH-1:0] a3_data_delayed_1;
wire [`DWIDTH-1:0] a3_data_delayed_2;
wire [`DWIDTH-1:0] a3_data_delayed_3;
wire [`DWIDTH-1:0] a4_data_delayed_1;
wire [`DWIDTH-1:0] a4_data_delayed_2;
wire [`DWIDTH-1:0] a4_data_delayed_3;
wire [`DWIDTH-1:0] a4_data_delayed_4;
wire [`DWIDTH-1:0] a5_data_delayed_1;
wire [`DWIDTH-1:0] a5_data_delayed_2;
wire [`DWIDTH-1:0] a5_data_delayed_3;
wire [`DWIDTH-1:0] a5_data_delayed_4;
wire [`DWIDTH-1:0] a5_data_delayed_5;
wire [`DWIDTH-1:0] a6_data_delayed_1;
wire [`DWIDTH-1:0] a6_data_delayed_2;
wire [`DWIDTH-1:0] a6_data_delayed_3;
wire [`DWIDTH-1:0] a6_data_delayed_4;
wire [`DWIDTH-1:0] a6_data_delayed_5;
wire [`DWIDTH-1:0] a6_data_delayed_6;
wire [`DWIDTH-1:0] a7_data_delayed_1;
wire [`DWIDTH-1:0] a7_data_delayed_2;
wire [`DWIDTH-1:0] a7_data_delayed_3;
wire [`DWIDTH-1:0] a7_data_delayed_4;
wire [`DWIDTH-1:0] a7_data_delayed_5;
wire [`DWIDTH-1:0] a7_data_delayed_6;
wire [`DWIDTH-1:0] a7_data_delayed_7;
wire [`DWIDTH-1:0] a8_data_delayed_1;
wire [`DWIDTH-1:0] a8_data_delayed_2;
wire [`DWIDTH-1:0] a8_data_delayed_3;
wire [`DWIDTH-1:0] a8_data_delayed_4;
wire [`DWIDTH-1:0] a8_data_delayed_5;
wire [`DWIDTH-1:0] a8_data_delayed_6;
wire [`DWIDTH-1:0] a8_data_delayed_7;
wire [`DWIDTH-1:0] a8_data_delayed_8;
wire [`DWIDTH-1:0] a9_data_delayed_1;
wire [`DWIDTH-1:0] a9_data_delayed_2;
wire [`DWIDTH-1:0] a9_data_delayed_3;
wire [`DWIDTH-1:0] a9_data_delayed_4;
wire [`DWIDTH-1:0] a9_data_delayed_5;
wire [`DWIDTH-1:0] a9_data_delayed_6;
wire [`DWIDTH-1:0] a9_data_delayed_7;
wire [`DWIDTH-1:0] a9_data_delayed_8;
wire [`DWIDTH-1:0] a9_data_delayed_9;
wire [`DWIDTH-1:0] a10_data_delayed_1;
wire [`DWIDTH-1:0] a10_data_delayed_2;
wire [`DWIDTH-1:0] a10_data_delayed_3;
wire [`DWIDTH-1:0] a10_data_delayed_4;
wire [`DWIDTH-1:0] a10_data_delayed_5;
wire [`DWIDTH-1:0] a10_data_delayed_6;
wire [`DWIDTH-1:0] a10_data_delayed_7;
wire [`DWIDTH-1:0] a10_data_delayed_8;
wire [`DWIDTH-1:0] a10_data_delayed_9;
wire [`DWIDTH-1:0] a10_data_delayed_10;
wire [`DWIDTH-1:0] a11_data_delayed_1;
wire [`DWIDTH-1:0] a11_data_delayed_2;
wire [`DWIDTH-1:0] a11_data_delayed_3;
wire [`DWIDTH-1:0] a11_data_delayed_4;
wire [`DWIDTH-1:0] a11_data_delayed_5;
wire [`DWIDTH-1:0] a11_data_delayed_6;
wire [`DWIDTH-1:0] a11_data_delayed_7;
wire [`DWIDTH-1:0] a11_data_delayed_8;
wire [`DWIDTH-1:0] a11_data_delayed_9;
wire [`DWIDTH-1:0] a11_data_delayed_10;
wire [`DWIDTH-1:0] a11_data_delayed_11;
wire [`DWIDTH-1:0] a12_data_delayed_1;
wire [`DWIDTH-1:0] a12_data_delayed_2;
wire [`DWIDTH-1:0] a12_data_delayed_3;
wire [`DWIDTH-1:0] a12_data_delayed_4;
wire [`DWIDTH-1:0] a12_data_delayed_5;
wire [`DWIDTH-1:0] a12_data_delayed_6;
wire [`DWIDTH-1:0] a12_data_delayed_7;
wire [`DWIDTH-1:0] a12_data_delayed_8;
wire [`DWIDTH-1:0] a12_data_delayed_9;
wire [`DWIDTH-1:0] a12_data_delayed_10;
wire [`DWIDTH-1:0] a12_data_delayed_11;
wire [`DWIDTH-1:0] a12_data_delayed_12;
wire [`DWIDTH-1:0] a13_data_delayed_1;
wire [`DWIDTH-1:0] a13_data_delayed_2;
wire [`DWIDTH-1:0] a13_data_delayed_3;
wire [`DWIDTH-1:0] a13_data_delayed_4;
wire [`DWIDTH-1:0] a13_data_delayed_5;
wire [`DWIDTH-1:0] a13_data_delayed_6;
wire [`DWIDTH-1:0] a13_data_delayed_7;
wire [`DWIDTH-1:0] a13_data_delayed_8;
wire [`DWIDTH-1:0] a13_data_delayed_9;
wire [`DWIDTH-1:0] a13_data_delayed_10;
wire [`DWIDTH-1:0] a13_data_delayed_11;
wire [`DWIDTH-1:0] a13_data_delayed_12;
wire [`DWIDTH-1:0] a13_data_delayed_13;
wire [`DWIDTH-1:0] a14_data_delayed_1;
wire [`DWIDTH-1:0] a14_data_delayed_2;
wire [`DWIDTH-1:0] a14_data_delayed_3;
wire [`DWIDTH-1:0] a14_data_delayed_4;
wire [`DWIDTH-1:0] a14_data_delayed_5;
wire [`DWIDTH-1:0] a14_data_delayed_6;
wire [`DWIDTH-1:0] a14_data_delayed_7;
wire [`DWIDTH-1:0] a14_data_delayed_8;
wire [`DWIDTH-1:0] a14_data_delayed_9;
wire [`DWIDTH-1:0] a14_data_delayed_10;
wire [`DWIDTH-1:0] a14_data_delayed_11;
wire [`DWIDTH-1:0] a14_data_delayed_12;
wire [`DWIDTH-1:0] a14_data_delayed_13;
wire [`DWIDTH-1:0] a14_data_delayed_14;
wire [`DWIDTH-1:0] a15_data_delayed_1;
wire [`DWIDTH-1:0] a15_data_delayed_2;
wire [`DWIDTH-1:0] a15_data_delayed_3;
wire [`DWIDTH-1:0] a15_data_delayed_4;
wire [`DWIDTH-1:0] a15_data_delayed_5;
wire [`DWIDTH-1:0] a15_data_delayed_6;
wire [`DWIDTH-1:0] a15_data_delayed_7;
wire [`DWIDTH-1:0] a15_data_delayed_8;
wire [`DWIDTH-1:0] a15_data_delayed_9;
wire [`DWIDTH-1:0] a15_data_delayed_10;
wire [`DWIDTH-1:0] a15_data_delayed_11;
wire [`DWIDTH-1:0] a15_data_delayed_12;
wire [`DWIDTH-1:0] a15_data_delayed_13;
wire [`DWIDTH-1:0] a15_data_delayed_14;
wire [`DWIDTH-1:0] a15_data_delayed_15;
wire [`DWIDTH-1:0] a16_data_delayed_1;
wire [`DWIDTH-1:0] a16_data_delayed_2;
wire [`DWIDTH-1:0] a16_data_delayed_3;
wire [`DWIDTH-1:0] a16_data_delayed_4;
wire [`DWIDTH-1:0] a16_data_delayed_5;
wire [`DWIDTH-1:0] a16_data_delayed_6;
wire [`DWIDTH-1:0] a16_data_delayed_7;
wire [`DWIDTH-1:0] a16_data_delayed_8;
wire [`DWIDTH-1:0] a16_data_delayed_9;
wire [`DWIDTH-1:0] a16_data_delayed_10;
wire [`DWIDTH-1:0] a16_data_delayed_11;
wire [`DWIDTH-1:0] a16_data_delayed_12;
wire [`DWIDTH-1:0] a16_data_delayed_13;
wire [`DWIDTH-1:0] a16_data_delayed_14;
wire [`DWIDTH-1:0] a16_data_delayed_15;
wire [`DWIDTH-1:0] a16_data_delayed_16;
wire [`DWIDTH-1:0] a17_data_delayed_1;
wire [`DWIDTH-1:0] a17_data_delayed_2;
wire [`DWIDTH-1:0] a17_data_delayed_3;
wire [`DWIDTH-1:0] a17_data_delayed_4;
wire [`DWIDTH-1:0] a17_data_delayed_5;
wire [`DWIDTH-1:0] a17_data_delayed_6;
wire [`DWIDTH-1:0] a17_data_delayed_7;
wire [`DWIDTH-1:0] a17_data_delayed_8;
wire [`DWIDTH-1:0] a17_data_delayed_9;
wire [`DWIDTH-1:0] a17_data_delayed_10;
wire [`DWIDTH-1:0] a17_data_delayed_11;
wire [`DWIDTH-1:0] a17_data_delayed_12;
wire [`DWIDTH-1:0] a17_data_delayed_13;
wire [`DWIDTH-1:0] a17_data_delayed_14;
wire [`DWIDTH-1:0] a17_data_delayed_15;
wire [`DWIDTH-1:0] a17_data_delayed_16;
wire [`DWIDTH-1:0] a17_data_delayed_17;
wire [`DWIDTH-1:0] a18_data_delayed_1;
wire [`DWIDTH-1:0] a18_data_delayed_2;
wire [`DWIDTH-1:0] a18_data_delayed_3;
wire [`DWIDTH-1:0] a18_data_delayed_4;
wire [`DWIDTH-1:0] a18_data_delayed_5;
wire [`DWIDTH-1:0] a18_data_delayed_6;
wire [`DWIDTH-1:0] a18_data_delayed_7;
wire [`DWIDTH-1:0] a18_data_delayed_8;
wire [`DWIDTH-1:0] a18_data_delayed_9;
wire [`DWIDTH-1:0] a18_data_delayed_10;
wire [`DWIDTH-1:0] a18_data_delayed_11;
wire [`DWIDTH-1:0] a18_data_delayed_12;
wire [`DWIDTH-1:0] a18_data_delayed_13;
wire [`DWIDTH-1:0] a18_data_delayed_14;
wire [`DWIDTH-1:0] a18_data_delayed_15;
wire [`DWIDTH-1:0] a18_data_delayed_16;
wire [`DWIDTH-1:0] a18_data_delayed_17;
wire [`DWIDTH-1:0] a18_data_delayed_18;
wire [`DWIDTH-1:0] a19_data_delayed_1;
wire [`DWIDTH-1:0] a19_data_delayed_2;
wire [`DWIDTH-1:0] a19_data_delayed_3;
wire [`DWIDTH-1:0] a19_data_delayed_4;
wire [`DWIDTH-1:0] a19_data_delayed_5;
wire [`DWIDTH-1:0] a19_data_delayed_6;
wire [`DWIDTH-1:0] a19_data_delayed_7;
wire [`DWIDTH-1:0] a19_data_delayed_8;
wire [`DWIDTH-1:0] a19_data_delayed_9;
wire [`DWIDTH-1:0] a19_data_delayed_10;
wire [`DWIDTH-1:0] a19_data_delayed_11;
wire [`DWIDTH-1:0] a19_data_delayed_12;
wire [`DWIDTH-1:0] a19_data_delayed_13;
wire [`DWIDTH-1:0] a19_data_delayed_14;
wire [`DWIDTH-1:0] a19_data_delayed_15;
wire [`DWIDTH-1:0] a19_data_delayed_16;
wire [`DWIDTH-1:0] a19_data_delayed_17;
wire [`DWIDTH-1:0] a19_data_delayed_18;
wire [`DWIDTH-1:0] a19_data_delayed_19;
wire [`DWIDTH-1:0] a20_data_delayed_1;
wire [`DWIDTH-1:0] a20_data_delayed_2;
wire [`DWIDTH-1:0] a20_data_delayed_3;
wire [`DWIDTH-1:0] a20_data_delayed_4;
wire [`DWIDTH-1:0] a20_data_delayed_5;
wire [`DWIDTH-1:0] a20_data_delayed_6;
wire [`DWIDTH-1:0] a20_data_delayed_7;
wire [`DWIDTH-1:0] a20_data_delayed_8;
wire [`DWIDTH-1:0] a20_data_delayed_9;
wire [`DWIDTH-1:0] a20_data_delayed_10;
wire [`DWIDTH-1:0] a20_data_delayed_11;
wire [`DWIDTH-1:0] a20_data_delayed_12;
wire [`DWIDTH-1:0] a20_data_delayed_13;
wire [`DWIDTH-1:0] a20_data_delayed_14;
wire [`DWIDTH-1:0] a20_data_delayed_15;
wire [`DWIDTH-1:0] a20_data_delayed_16;
wire [`DWIDTH-1:0] a20_data_delayed_17;
wire [`DWIDTH-1:0] a20_data_delayed_18;
wire [`DWIDTH-1:0] a20_data_delayed_19;
wire [`DWIDTH-1:0] a20_data_delayed_20;
wire [`DWIDTH-1:0] a21_data_delayed_1;
wire [`DWIDTH-1:0] a21_data_delayed_2;
wire [`DWIDTH-1:0] a21_data_delayed_3;
wire [`DWIDTH-1:0] a21_data_delayed_4;
wire [`DWIDTH-1:0] a21_data_delayed_5;
wire [`DWIDTH-1:0] a21_data_delayed_6;
wire [`DWIDTH-1:0] a21_data_delayed_7;
wire [`DWIDTH-1:0] a21_data_delayed_8;
wire [`DWIDTH-1:0] a21_data_delayed_9;
wire [`DWIDTH-1:0] a21_data_delayed_10;
wire [`DWIDTH-1:0] a21_data_delayed_11;
wire [`DWIDTH-1:0] a21_data_delayed_12;
wire [`DWIDTH-1:0] a21_data_delayed_13;
wire [`DWIDTH-1:0] a21_data_delayed_14;
wire [`DWIDTH-1:0] a21_data_delayed_15;
wire [`DWIDTH-1:0] a21_data_delayed_16;
wire [`DWIDTH-1:0] a21_data_delayed_17;
wire [`DWIDTH-1:0] a21_data_delayed_18;
wire [`DWIDTH-1:0] a21_data_delayed_19;
wire [`DWIDTH-1:0] a21_data_delayed_20;
wire [`DWIDTH-1:0] a21_data_delayed_21;
wire [`DWIDTH-1:0] a22_data_delayed_1;
wire [`DWIDTH-1:0] a22_data_delayed_2;
wire [`DWIDTH-1:0] a22_data_delayed_3;
wire [`DWIDTH-1:0] a22_data_delayed_4;
wire [`DWIDTH-1:0] a22_data_delayed_5;
wire [`DWIDTH-1:0] a22_data_delayed_6;
wire [`DWIDTH-1:0] a22_data_delayed_7;
wire [`DWIDTH-1:0] a22_data_delayed_8;
wire [`DWIDTH-1:0] a22_data_delayed_9;
wire [`DWIDTH-1:0] a22_data_delayed_10;
wire [`DWIDTH-1:0] a22_data_delayed_11;
wire [`DWIDTH-1:0] a22_data_delayed_12;
wire [`DWIDTH-1:0] a22_data_delayed_13;
wire [`DWIDTH-1:0] a22_data_delayed_14;
wire [`DWIDTH-1:0] a22_data_delayed_15;
wire [`DWIDTH-1:0] a22_data_delayed_16;
wire [`DWIDTH-1:0] a22_data_delayed_17;
wire [`DWIDTH-1:0] a22_data_delayed_18;
wire [`DWIDTH-1:0] a22_data_delayed_19;
wire [`DWIDTH-1:0] a22_data_delayed_20;
wire [`DWIDTH-1:0] a22_data_delayed_21;
wire [`DWIDTH-1:0] a22_data_delayed_22;
wire [`DWIDTH-1:0] a23_data_delayed_1;
wire [`DWIDTH-1:0] a23_data_delayed_2;
wire [`DWIDTH-1:0] a23_data_delayed_3;
wire [`DWIDTH-1:0] a23_data_delayed_4;
wire [`DWIDTH-1:0] a23_data_delayed_5;
wire [`DWIDTH-1:0] a23_data_delayed_6;
wire [`DWIDTH-1:0] a23_data_delayed_7;
wire [`DWIDTH-1:0] a23_data_delayed_8;
wire [`DWIDTH-1:0] a23_data_delayed_9;
wire [`DWIDTH-1:0] a23_data_delayed_10;
wire [`DWIDTH-1:0] a23_data_delayed_11;
wire [`DWIDTH-1:0] a23_data_delayed_12;
wire [`DWIDTH-1:0] a23_data_delayed_13;
wire [`DWIDTH-1:0] a23_data_delayed_14;
wire [`DWIDTH-1:0] a23_data_delayed_15;
wire [`DWIDTH-1:0] a23_data_delayed_16;
wire [`DWIDTH-1:0] a23_data_delayed_17;
wire [`DWIDTH-1:0] a23_data_delayed_18;
wire [`DWIDTH-1:0] a23_data_delayed_19;
wire [`DWIDTH-1:0] a23_data_delayed_20;
wire [`DWIDTH-1:0] a23_data_delayed_21;
wire [`DWIDTH-1:0] a23_data_delayed_22;
wire [`DWIDTH-1:0] a23_data_delayed_23;
wire [`DWIDTH-1:0] a24_data_delayed_1;
wire [`DWIDTH-1:0] a24_data_delayed_2;
wire [`DWIDTH-1:0] a24_data_delayed_3;
wire [`DWIDTH-1:0] a24_data_delayed_4;
wire [`DWIDTH-1:0] a24_data_delayed_5;
wire [`DWIDTH-1:0] a24_data_delayed_6;
wire [`DWIDTH-1:0] a24_data_delayed_7;
wire [`DWIDTH-1:0] a24_data_delayed_8;
wire [`DWIDTH-1:0] a24_data_delayed_9;
wire [`DWIDTH-1:0] a24_data_delayed_10;
wire [`DWIDTH-1:0] a24_data_delayed_11;
wire [`DWIDTH-1:0] a24_data_delayed_12;
wire [`DWIDTH-1:0] a24_data_delayed_13;
wire [`DWIDTH-1:0] a24_data_delayed_14;
wire [`DWIDTH-1:0] a24_data_delayed_15;
wire [`DWIDTH-1:0] a24_data_delayed_16;
wire [`DWIDTH-1:0] a24_data_delayed_17;
wire [`DWIDTH-1:0] a24_data_delayed_18;
wire [`DWIDTH-1:0] a24_data_delayed_19;
wire [`DWIDTH-1:0] a24_data_delayed_20;
wire [`DWIDTH-1:0] a24_data_delayed_21;
wire [`DWIDTH-1:0] a24_data_delayed_22;
wire [`DWIDTH-1:0] a24_data_delayed_23;
wire [`DWIDTH-1:0] a24_data_delayed_24;
wire [`DWIDTH-1:0] a25_data_delayed_1;
wire [`DWIDTH-1:0] a25_data_delayed_2;
wire [`DWIDTH-1:0] a25_data_delayed_3;
wire [`DWIDTH-1:0] a25_data_delayed_4;
wire [`DWIDTH-1:0] a25_data_delayed_5;
wire [`DWIDTH-1:0] a25_data_delayed_6;
wire [`DWIDTH-1:0] a25_data_delayed_7;
wire [`DWIDTH-1:0] a25_data_delayed_8;
wire [`DWIDTH-1:0] a25_data_delayed_9;
wire [`DWIDTH-1:0] a25_data_delayed_10;
wire [`DWIDTH-1:0] a25_data_delayed_11;
wire [`DWIDTH-1:0] a25_data_delayed_12;
wire [`DWIDTH-1:0] a25_data_delayed_13;
wire [`DWIDTH-1:0] a25_data_delayed_14;
wire [`DWIDTH-1:0] a25_data_delayed_15;
wire [`DWIDTH-1:0] a25_data_delayed_16;
wire [`DWIDTH-1:0] a25_data_delayed_17;
wire [`DWIDTH-1:0] a25_data_delayed_18;
wire [`DWIDTH-1:0] a25_data_delayed_19;
wire [`DWIDTH-1:0] a25_data_delayed_20;
wire [`DWIDTH-1:0] a25_data_delayed_21;
wire [`DWIDTH-1:0] a25_data_delayed_22;
wire [`DWIDTH-1:0] a25_data_delayed_23;
wire [`DWIDTH-1:0] a25_data_delayed_24;
wire [`DWIDTH-1:0] a25_data_delayed_25;
wire [`DWIDTH-1:0] a26_data_delayed_1;
wire [`DWIDTH-1:0] a26_data_delayed_2;
wire [`DWIDTH-1:0] a26_data_delayed_3;
wire [`DWIDTH-1:0] a26_data_delayed_4;
wire [`DWIDTH-1:0] a26_data_delayed_5;
wire [`DWIDTH-1:0] a26_data_delayed_6;
wire [`DWIDTH-1:0] a26_data_delayed_7;
wire [`DWIDTH-1:0] a26_data_delayed_8;
wire [`DWIDTH-1:0] a26_data_delayed_9;
wire [`DWIDTH-1:0] a26_data_delayed_10;
wire [`DWIDTH-1:0] a26_data_delayed_11;
wire [`DWIDTH-1:0] a26_data_delayed_12;
wire [`DWIDTH-1:0] a26_data_delayed_13;
wire [`DWIDTH-1:0] a26_data_delayed_14;
wire [`DWIDTH-1:0] a26_data_delayed_15;
wire [`DWIDTH-1:0] a26_data_delayed_16;
wire [`DWIDTH-1:0] a26_data_delayed_17;
wire [`DWIDTH-1:0] a26_data_delayed_18;
wire [`DWIDTH-1:0] a26_data_delayed_19;
wire [`DWIDTH-1:0] a26_data_delayed_20;
wire [`DWIDTH-1:0] a26_data_delayed_21;
wire [`DWIDTH-1:0] a26_data_delayed_22;
wire [`DWIDTH-1:0] a26_data_delayed_23;
wire [`DWIDTH-1:0] a26_data_delayed_24;
wire [`DWIDTH-1:0] a26_data_delayed_25;
wire [`DWIDTH-1:0] a26_data_delayed_26;
wire [`DWIDTH-1:0] a27_data_delayed_1;
wire [`DWIDTH-1:0] a27_data_delayed_2;
wire [`DWIDTH-1:0] a27_data_delayed_3;
wire [`DWIDTH-1:0] a27_data_delayed_4;
wire [`DWIDTH-1:0] a27_data_delayed_5;
wire [`DWIDTH-1:0] a27_data_delayed_6;
wire [`DWIDTH-1:0] a27_data_delayed_7;
wire [`DWIDTH-1:0] a27_data_delayed_8;
wire [`DWIDTH-1:0] a27_data_delayed_9;
wire [`DWIDTH-1:0] a27_data_delayed_10;
wire [`DWIDTH-1:0] a27_data_delayed_11;
wire [`DWIDTH-1:0] a27_data_delayed_12;
wire [`DWIDTH-1:0] a27_data_delayed_13;
wire [`DWIDTH-1:0] a27_data_delayed_14;
wire [`DWIDTH-1:0] a27_data_delayed_15;
wire [`DWIDTH-1:0] a27_data_delayed_16;
wire [`DWIDTH-1:0] a27_data_delayed_17;
wire [`DWIDTH-1:0] a27_data_delayed_18;
wire [`DWIDTH-1:0] a27_data_delayed_19;
wire [`DWIDTH-1:0] a27_data_delayed_20;
wire [`DWIDTH-1:0] a27_data_delayed_21;
wire [`DWIDTH-1:0] a27_data_delayed_22;
wire [`DWIDTH-1:0] a27_data_delayed_23;
wire [`DWIDTH-1:0] a27_data_delayed_24;
wire [`DWIDTH-1:0] a27_data_delayed_25;
wire [`DWIDTH-1:0] a27_data_delayed_26;
wire [`DWIDTH-1:0] a27_data_delayed_27;
wire [`DWIDTH-1:0] a28_data_delayed_1;
wire [`DWIDTH-1:0] a28_data_delayed_2;
wire [`DWIDTH-1:0] a28_data_delayed_3;
wire [`DWIDTH-1:0] a28_data_delayed_4;
wire [`DWIDTH-1:0] a28_data_delayed_5;
wire [`DWIDTH-1:0] a28_data_delayed_6;
wire [`DWIDTH-1:0] a28_data_delayed_7;
wire [`DWIDTH-1:0] a28_data_delayed_8;
wire [`DWIDTH-1:0] a28_data_delayed_9;
wire [`DWIDTH-1:0] a28_data_delayed_10;
wire [`DWIDTH-1:0] a28_data_delayed_11;
wire [`DWIDTH-1:0] a28_data_delayed_12;
wire [`DWIDTH-1:0] a28_data_delayed_13;
wire [`DWIDTH-1:0] a28_data_delayed_14;
wire [`DWIDTH-1:0] a28_data_delayed_15;
wire [`DWIDTH-1:0] a28_data_delayed_16;
wire [`DWIDTH-1:0] a28_data_delayed_17;
wire [`DWIDTH-1:0] a28_data_delayed_18;
wire [`DWIDTH-1:0] a28_data_delayed_19;
wire [`DWIDTH-1:0] a28_data_delayed_20;
wire [`DWIDTH-1:0] a28_data_delayed_21;
wire [`DWIDTH-1:0] a28_data_delayed_22;
wire [`DWIDTH-1:0] a28_data_delayed_23;
wire [`DWIDTH-1:0] a28_data_delayed_24;
wire [`DWIDTH-1:0] a28_data_delayed_25;
wire [`DWIDTH-1:0] a28_data_delayed_26;
wire [`DWIDTH-1:0] a28_data_delayed_27;
wire [`DWIDTH-1:0] a28_data_delayed_28;
wire [`DWIDTH-1:0] a29_data_delayed_1;
wire [`DWIDTH-1:0] a29_data_delayed_2;
wire [`DWIDTH-1:0] a29_data_delayed_3;
wire [`DWIDTH-1:0] a29_data_delayed_4;
wire [`DWIDTH-1:0] a29_data_delayed_5;
wire [`DWIDTH-1:0] a29_data_delayed_6;
wire [`DWIDTH-1:0] a29_data_delayed_7;
wire [`DWIDTH-1:0] a29_data_delayed_8;
wire [`DWIDTH-1:0] a29_data_delayed_9;
wire [`DWIDTH-1:0] a29_data_delayed_10;
wire [`DWIDTH-1:0] a29_data_delayed_11;
wire [`DWIDTH-1:0] a29_data_delayed_12;
wire [`DWIDTH-1:0] a29_data_delayed_13;
wire [`DWIDTH-1:0] a29_data_delayed_14;
wire [`DWIDTH-1:0] a29_data_delayed_15;
wire [`DWIDTH-1:0] a29_data_delayed_16;
wire [`DWIDTH-1:0] a29_data_delayed_17;
wire [`DWIDTH-1:0] a29_data_delayed_18;
wire [`DWIDTH-1:0] a29_data_delayed_19;
wire [`DWIDTH-1:0] a29_data_delayed_20;
wire [`DWIDTH-1:0] a29_data_delayed_21;
wire [`DWIDTH-1:0] a29_data_delayed_22;
wire [`DWIDTH-1:0] a29_data_delayed_23;
wire [`DWIDTH-1:0] a29_data_delayed_24;
wire [`DWIDTH-1:0] a29_data_delayed_25;
wire [`DWIDTH-1:0] a29_data_delayed_26;
wire [`DWIDTH-1:0] a29_data_delayed_27;
wire [`DWIDTH-1:0] a29_data_delayed_28;
wire [`DWIDTH-1:0] a29_data_delayed_29;
wire [`DWIDTH-1:0] a30_data_delayed_1;
wire [`DWIDTH-1:0] a30_data_delayed_2;
wire [`DWIDTH-1:0] a30_data_delayed_3;
wire [`DWIDTH-1:0] a30_data_delayed_4;
wire [`DWIDTH-1:0] a30_data_delayed_5;
wire [`DWIDTH-1:0] a30_data_delayed_6;
wire [`DWIDTH-1:0] a30_data_delayed_7;
wire [`DWIDTH-1:0] a30_data_delayed_8;
wire [`DWIDTH-1:0] a30_data_delayed_9;
wire [`DWIDTH-1:0] a30_data_delayed_10;
wire [`DWIDTH-1:0] a30_data_delayed_11;
wire [`DWIDTH-1:0] a30_data_delayed_12;
wire [`DWIDTH-1:0] a30_data_delayed_13;
wire [`DWIDTH-1:0] a30_data_delayed_14;
wire [`DWIDTH-1:0] a30_data_delayed_15;
wire [`DWIDTH-1:0] a30_data_delayed_16;
wire [`DWIDTH-1:0] a30_data_delayed_17;
wire [`DWIDTH-1:0] a30_data_delayed_18;
wire [`DWIDTH-1:0] a30_data_delayed_19;
wire [`DWIDTH-1:0] a30_data_delayed_20;
wire [`DWIDTH-1:0] a30_data_delayed_21;
wire [`DWIDTH-1:0] a30_data_delayed_22;
wire [`DWIDTH-1:0] a30_data_delayed_23;
wire [`DWIDTH-1:0] a30_data_delayed_24;
wire [`DWIDTH-1:0] a30_data_delayed_25;
wire [`DWIDTH-1:0] a30_data_delayed_26;
wire [`DWIDTH-1:0] a30_data_delayed_27;
wire [`DWIDTH-1:0] a30_data_delayed_28;
wire [`DWIDTH-1:0] a30_data_delayed_29;
wire [`DWIDTH-1:0] a30_data_delayed_30;
wire [`DWIDTH-1:0] a31_data_delayed_1;
wire [`DWIDTH-1:0] a31_data_delayed_2;
wire [`DWIDTH-1:0] a31_data_delayed_3;
wire [`DWIDTH-1:0] a31_data_delayed_4;
wire [`DWIDTH-1:0] a31_data_delayed_5;
wire [`DWIDTH-1:0] a31_data_delayed_6;
wire [`DWIDTH-1:0] a31_data_delayed_7;
wire [`DWIDTH-1:0] a31_data_delayed_8;
wire [`DWIDTH-1:0] a31_data_delayed_9;
wire [`DWIDTH-1:0] a31_data_delayed_10;
wire [`DWIDTH-1:0] a31_data_delayed_11;
wire [`DWIDTH-1:0] a31_data_delayed_12;
wire [`DWIDTH-1:0] a31_data_delayed_13;
wire [`DWIDTH-1:0] a31_data_delayed_14;
wire [`DWIDTH-1:0] a31_data_delayed_15;
wire [`DWIDTH-1:0] a31_data_delayed_16;
wire [`DWIDTH-1:0] a31_data_delayed_17;
wire [`DWIDTH-1:0] a31_data_delayed_18;
wire [`DWIDTH-1:0] a31_data_delayed_19;
wire [`DWIDTH-1:0] a31_data_delayed_20;
wire [`DWIDTH-1:0] a31_data_delayed_21;
wire [`DWIDTH-1:0] a31_data_delayed_22;
wire [`DWIDTH-1:0] a31_data_delayed_23;
wire [`DWIDTH-1:0] a31_data_delayed_24;
wire [`DWIDTH-1:0] a31_data_delayed_25;
wire [`DWIDTH-1:0] a31_data_delayed_26;
wire [`DWIDTH-1:0] a31_data_delayed_27;
wire [`DWIDTH-1:0] a31_data_delayed_28;
wire [`DWIDTH-1:0] a31_data_delayed_29;
wire [`DWIDTH-1:0] a31_data_delayed_30;
wire [`DWIDTH-1:0] a31_data_delayed_31;
wire [`DWIDTH-1:0] b1_data_delayed_1;
wire [`DWIDTH-1:0] b2_data_delayed_1;
wire [`DWIDTH-1:0] b2_data_delayed_2;
wire [`DWIDTH-1:0] b3_data_delayed_1;
wire [`DWIDTH-1:0] b3_data_delayed_2;
wire [`DWIDTH-1:0] b3_data_delayed_3;
wire [`DWIDTH-1:0] b4_data_delayed_1;
wire [`DWIDTH-1:0] b4_data_delayed_2;
wire [`DWIDTH-1:0] b4_data_delayed_3;
wire [`DWIDTH-1:0] b4_data_delayed_4;
wire [`DWIDTH-1:0] b5_data_delayed_1;
wire [`DWIDTH-1:0] b5_data_delayed_2;
wire [`DWIDTH-1:0] b5_data_delayed_3;
wire [`DWIDTH-1:0] b5_data_delayed_4;
wire [`DWIDTH-1:0] b5_data_delayed_5;
wire [`DWIDTH-1:0] b6_data_delayed_1;
wire [`DWIDTH-1:0] b6_data_delayed_2;
wire [`DWIDTH-1:0] b6_data_delayed_3;
wire [`DWIDTH-1:0] b6_data_delayed_4;
wire [`DWIDTH-1:0] b6_data_delayed_5;
wire [`DWIDTH-1:0] b6_data_delayed_6;
wire [`DWIDTH-1:0] b7_data_delayed_1;
wire [`DWIDTH-1:0] b7_data_delayed_2;
wire [`DWIDTH-1:0] b7_data_delayed_3;
wire [`DWIDTH-1:0] b7_data_delayed_4;
wire [`DWIDTH-1:0] b7_data_delayed_5;
wire [`DWIDTH-1:0] b7_data_delayed_6;
wire [`DWIDTH-1:0] b7_data_delayed_7;
wire [`DWIDTH-1:0] b8_data_delayed_1;
wire [`DWIDTH-1:0] b8_data_delayed_2;
wire [`DWIDTH-1:0] b8_data_delayed_3;
wire [`DWIDTH-1:0] b8_data_delayed_4;
wire [`DWIDTH-1:0] b8_data_delayed_5;
wire [`DWIDTH-1:0] b8_data_delayed_6;
wire [`DWIDTH-1:0] b8_data_delayed_7;
wire [`DWIDTH-1:0] b8_data_delayed_8;
wire [`DWIDTH-1:0] b9_data_delayed_1;
wire [`DWIDTH-1:0] b9_data_delayed_2;
wire [`DWIDTH-1:0] b9_data_delayed_3;
wire [`DWIDTH-1:0] b9_data_delayed_4;
wire [`DWIDTH-1:0] b9_data_delayed_5;
wire [`DWIDTH-1:0] b9_data_delayed_6;
wire [`DWIDTH-1:0] b9_data_delayed_7;
wire [`DWIDTH-1:0] b9_data_delayed_8;
wire [`DWIDTH-1:0] b9_data_delayed_9;
wire [`DWIDTH-1:0] b10_data_delayed_1;
wire [`DWIDTH-1:0] b10_data_delayed_2;
wire [`DWIDTH-1:0] b10_data_delayed_3;
wire [`DWIDTH-1:0] b10_data_delayed_4;
wire [`DWIDTH-1:0] b10_data_delayed_5;
wire [`DWIDTH-1:0] b10_data_delayed_6;
wire [`DWIDTH-1:0] b10_data_delayed_7;
wire [`DWIDTH-1:0] b10_data_delayed_8;
wire [`DWIDTH-1:0] b10_data_delayed_9;
wire [`DWIDTH-1:0] b10_data_delayed_10;
wire [`DWIDTH-1:0] b11_data_delayed_1;
wire [`DWIDTH-1:0] b11_data_delayed_2;
wire [`DWIDTH-1:0] b11_data_delayed_3;
wire [`DWIDTH-1:0] b11_data_delayed_4;
wire [`DWIDTH-1:0] b11_data_delayed_5;
wire [`DWIDTH-1:0] b11_data_delayed_6;
wire [`DWIDTH-1:0] b11_data_delayed_7;
wire [`DWIDTH-1:0] b11_data_delayed_8;
wire [`DWIDTH-1:0] b11_data_delayed_9;
wire [`DWIDTH-1:0] b11_data_delayed_10;
wire [`DWIDTH-1:0] b11_data_delayed_11;
wire [`DWIDTH-1:0] b12_data_delayed_1;
wire [`DWIDTH-1:0] b12_data_delayed_2;
wire [`DWIDTH-1:0] b12_data_delayed_3;
wire [`DWIDTH-1:0] b12_data_delayed_4;
wire [`DWIDTH-1:0] b12_data_delayed_5;
wire [`DWIDTH-1:0] b12_data_delayed_6;
wire [`DWIDTH-1:0] b12_data_delayed_7;
wire [`DWIDTH-1:0] b12_data_delayed_8;
wire [`DWIDTH-1:0] b12_data_delayed_9;
wire [`DWIDTH-1:0] b12_data_delayed_10;
wire [`DWIDTH-1:0] b12_data_delayed_11;
wire [`DWIDTH-1:0] b12_data_delayed_12;
wire [`DWIDTH-1:0] b13_data_delayed_1;
wire [`DWIDTH-1:0] b13_data_delayed_2;
wire [`DWIDTH-1:0] b13_data_delayed_3;
wire [`DWIDTH-1:0] b13_data_delayed_4;
wire [`DWIDTH-1:0] b13_data_delayed_5;
wire [`DWIDTH-1:0] b13_data_delayed_6;
wire [`DWIDTH-1:0] b13_data_delayed_7;
wire [`DWIDTH-1:0] b13_data_delayed_8;
wire [`DWIDTH-1:0] b13_data_delayed_9;
wire [`DWIDTH-1:0] b13_data_delayed_10;
wire [`DWIDTH-1:0] b13_data_delayed_11;
wire [`DWIDTH-1:0] b13_data_delayed_12;
wire [`DWIDTH-1:0] b13_data_delayed_13;
wire [`DWIDTH-1:0] b14_data_delayed_1;
wire [`DWIDTH-1:0] b14_data_delayed_2;
wire [`DWIDTH-1:0] b14_data_delayed_3;
wire [`DWIDTH-1:0] b14_data_delayed_4;
wire [`DWIDTH-1:0] b14_data_delayed_5;
wire [`DWIDTH-1:0] b14_data_delayed_6;
wire [`DWIDTH-1:0] b14_data_delayed_7;
wire [`DWIDTH-1:0] b14_data_delayed_8;
wire [`DWIDTH-1:0] b14_data_delayed_9;
wire [`DWIDTH-1:0] b14_data_delayed_10;
wire [`DWIDTH-1:0] b14_data_delayed_11;
wire [`DWIDTH-1:0] b14_data_delayed_12;
wire [`DWIDTH-1:0] b14_data_delayed_13;
wire [`DWIDTH-1:0] b14_data_delayed_14;
wire [`DWIDTH-1:0] b15_data_delayed_1;
wire [`DWIDTH-1:0] b15_data_delayed_2;
wire [`DWIDTH-1:0] b15_data_delayed_3;
wire [`DWIDTH-1:0] b15_data_delayed_4;
wire [`DWIDTH-1:0] b15_data_delayed_5;
wire [`DWIDTH-1:0] b15_data_delayed_6;
wire [`DWIDTH-1:0] b15_data_delayed_7;
wire [`DWIDTH-1:0] b15_data_delayed_8;
wire [`DWIDTH-1:0] b15_data_delayed_9;
wire [`DWIDTH-1:0] b15_data_delayed_10;
wire [`DWIDTH-1:0] b15_data_delayed_11;
wire [`DWIDTH-1:0] b15_data_delayed_12;
wire [`DWIDTH-1:0] b15_data_delayed_13;
wire [`DWIDTH-1:0] b15_data_delayed_14;
wire [`DWIDTH-1:0] b15_data_delayed_15;
wire [`DWIDTH-1:0] b16_data_delayed_1;
wire [`DWIDTH-1:0] b16_data_delayed_2;
wire [`DWIDTH-1:0] b16_data_delayed_3;
wire [`DWIDTH-1:0] b16_data_delayed_4;
wire [`DWIDTH-1:0] b16_data_delayed_5;
wire [`DWIDTH-1:0] b16_data_delayed_6;
wire [`DWIDTH-1:0] b16_data_delayed_7;
wire [`DWIDTH-1:0] b16_data_delayed_8;
wire [`DWIDTH-1:0] b16_data_delayed_9;
wire [`DWIDTH-1:0] b16_data_delayed_10;
wire [`DWIDTH-1:0] b16_data_delayed_11;
wire [`DWIDTH-1:0] b16_data_delayed_12;
wire [`DWIDTH-1:0] b16_data_delayed_13;
wire [`DWIDTH-1:0] b16_data_delayed_14;
wire [`DWIDTH-1:0] b16_data_delayed_15;
wire [`DWIDTH-1:0] b16_data_delayed_16;
wire [`DWIDTH-1:0] b17_data_delayed_1;
wire [`DWIDTH-1:0] b17_data_delayed_2;
wire [`DWIDTH-1:0] b17_data_delayed_3;
wire [`DWIDTH-1:0] b17_data_delayed_4;
wire [`DWIDTH-1:0] b17_data_delayed_5;
wire [`DWIDTH-1:0] b17_data_delayed_6;
wire [`DWIDTH-1:0] b17_data_delayed_7;
wire [`DWIDTH-1:0] b17_data_delayed_8;
wire [`DWIDTH-1:0] b17_data_delayed_9;
wire [`DWIDTH-1:0] b17_data_delayed_10;
wire [`DWIDTH-1:0] b17_data_delayed_11;
wire [`DWIDTH-1:0] b17_data_delayed_12;
wire [`DWIDTH-1:0] b17_data_delayed_13;
wire [`DWIDTH-1:0] b17_data_delayed_14;
wire [`DWIDTH-1:0] b17_data_delayed_15;
wire [`DWIDTH-1:0] b17_data_delayed_16;
wire [`DWIDTH-1:0] b17_data_delayed_17;
wire [`DWIDTH-1:0] b18_data_delayed_1;
wire [`DWIDTH-1:0] b18_data_delayed_2;
wire [`DWIDTH-1:0] b18_data_delayed_3;
wire [`DWIDTH-1:0] b18_data_delayed_4;
wire [`DWIDTH-1:0] b18_data_delayed_5;
wire [`DWIDTH-1:0] b18_data_delayed_6;
wire [`DWIDTH-1:0] b18_data_delayed_7;
wire [`DWIDTH-1:0] b18_data_delayed_8;
wire [`DWIDTH-1:0] b18_data_delayed_9;
wire [`DWIDTH-1:0] b18_data_delayed_10;
wire [`DWIDTH-1:0] b18_data_delayed_11;
wire [`DWIDTH-1:0] b18_data_delayed_12;
wire [`DWIDTH-1:0] b18_data_delayed_13;
wire [`DWIDTH-1:0] b18_data_delayed_14;
wire [`DWIDTH-1:0] b18_data_delayed_15;
wire [`DWIDTH-1:0] b18_data_delayed_16;
wire [`DWIDTH-1:0] b18_data_delayed_17;
wire [`DWIDTH-1:0] b18_data_delayed_18;
wire [`DWIDTH-1:0] b19_data_delayed_1;
wire [`DWIDTH-1:0] b19_data_delayed_2;
wire [`DWIDTH-1:0] b19_data_delayed_3;
wire [`DWIDTH-1:0] b19_data_delayed_4;
wire [`DWIDTH-1:0] b19_data_delayed_5;
wire [`DWIDTH-1:0] b19_data_delayed_6;
wire [`DWIDTH-1:0] b19_data_delayed_7;
wire [`DWIDTH-1:0] b19_data_delayed_8;
wire [`DWIDTH-1:0] b19_data_delayed_9;
wire [`DWIDTH-1:0] b19_data_delayed_10;
wire [`DWIDTH-1:0] b19_data_delayed_11;
wire [`DWIDTH-1:0] b19_data_delayed_12;
wire [`DWIDTH-1:0] b19_data_delayed_13;
wire [`DWIDTH-1:0] b19_data_delayed_14;
wire [`DWIDTH-1:0] b19_data_delayed_15;
wire [`DWIDTH-1:0] b19_data_delayed_16;
wire [`DWIDTH-1:0] b19_data_delayed_17;
wire [`DWIDTH-1:0] b19_data_delayed_18;
wire [`DWIDTH-1:0] b19_data_delayed_19;
wire [`DWIDTH-1:0] b20_data_delayed_1;
wire [`DWIDTH-1:0] b20_data_delayed_2;
wire [`DWIDTH-1:0] b20_data_delayed_3;
wire [`DWIDTH-1:0] b20_data_delayed_4;
wire [`DWIDTH-1:0] b20_data_delayed_5;
wire [`DWIDTH-1:0] b20_data_delayed_6;
wire [`DWIDTH-1:0] b20_data_delayed_7;
wire [`DWIDTH-1:0] b20_data_delayed_8;
wire [`DWIDTH-1:0] b20_data_delayed_9;
wire [`DWIDTH-1:0] b20_data_delayed_10;
wire [`DWIDTH-1:0] b20_data_delayed_11;
wire [`DWIDTH-1:0] b20_data_delayed_12;
wire [`DWIDTH-1:0] b20_data_delayed_13;
wire [`DWIDTH-1:0] b20_data_delayed_14;
wire [`DWIDTH-1:0] b20_data_delayed_15;
wire [`DWIDTH-1:0] b20_data_delayed_16;
wire [`DWIDTH-1:0] b20_data_delayed_17;
wire [`DWIDTH-1:0] b20_data_delayed_18;
wire [`DWIDTH-1:0] b20_data_delayed_19;
wire [`DWIDTH-1:0] b20_data_delayed_20;
wire [`DWIDTH-1:0] b21_data_delayed_1;
wire [`DWIDTH-1:0] b21_data_delayed_2;
wire [`DWIDTH-1:0] b21_data_delayed_3;
wire [`DWIDTH-1:0] b21_data_delayed_4;
wire [`DWIDTH-1:0] b21_data_delayed_5;
wire [`DWIDTH-1:0] b21_data_delayed_6;
wire [`DWIDTH-1:0] b21_data_delayed_7;
wire [`DWIDTH-1:0] b21_data_delayed_8;
wire [`DWIDTH-1:0] b21_data_delayed_9;
wire [`DWIDTH-1:0] b21_data_delayed_10;
wire [`DWIDTH-1:0] b21_data_delayed_11;
wire [`DWIDTH-1:0] b21_data_delayed_12;
wire [`DWIDTH-1:0] b21_data_delayed_13;
wire [`DWIDTH-1:0] b21_data_delayed_14;
wire [`DWIDTH-1:0] b21_data_delayed_15;
wire [`DWIDTH-1:0] b21_data_delayed_16;
wire [`DWIDTH-1:0] b21_data_delayed_17;
wire [`DWIDTH-1:0] b21_data_delayed_18;
wire [`DWIDTH-1:0] b21_data_delayed_19;
wire [`DWIDTH-1:0] b21_data_delayed_20;
wire [`DWIDTH-1:0] b21_data_delayed_21;
wire [`DWIDTH-1:0] b22_data_delayed_1;
wire [`DWIDTH-1:0] b22_data_delayed_2;
wire [`DWIDTH-1:0] b22_data_delayed_3;
wire [`DWIDTH-1:0] b22_data_delayed_4;
wire [`DWIDTH-1:0] b22_data_delayed_5;
wire [`DWIDTH-1:0] b22_data_delayed_6;
wire [`DWIDTH-1:0] b22_data_delayed_7;
wire [`DWIDTH-1:0] b22_data_delayed_8;
wire [`DWIDTH-1:0] b22_data_delayed_9;
wire [`DWIDTH-1:0] b22_data_delayed_10;
wire [`DWIDTH-1:0] b22_data_delayed_11;
wire [`DWIDTH-1:0] b22_data_delayed_12;
wire [`DWIDTH-1:0] b22_data_delayed_13;
wire [`DWIDTH-1:0] b22_data_delayed_14;
wire [`DWIDTH-1:0] b22_data_delayed_15;
wire [`DWIDTH-1:0] b22_data_delayed_16;
wire [`DWIDTH-1:0] b22_data_delayed_17;
wire [`DWIDTH-1:0] b22_data_delayed_18;
wire [`DWIDTH-1:0] b22_data_delayed_19;
wire [`DWIDTH-1:0] b22_data_delayed_20;
wire [`DWIDTH-1:0] b22_data_delayed_21;
wire [`DWIDTH-1:0] b22_data_delayed_22;
wire [`DWIDTH-1:0] b23_data_delayed_1;
wire [`DWIDTH-1:0] b23_data_delayed_2;
wire [`DWIDTH-1:0] b23_data_delayed_3;
wire [`DWIDTH-1:0] b23_data_delayed_4;
wire [`DWIDTH-1:0] b23_data_delayed_5;
wire [`DWIDTH-1:0] b23_data_delayed_6;
wire [`DWIDTH-1:0] b23_data_delayed_7;
wire [`DWIDTH-1:0] b23_data_delayed_8;
wire [`DWIDTH-1:0] b23_data_delayed_9;
wire [`DWIDTH-1:0] b23_data_delayed_10;
wire [`DWIDTH-1:0] b23_data_delayed_11;
wire [`DWIDTH-1:0] b23_data_delayed_12;
wire [`DWIDTH-1:0] b23_data_delayed_13;
wire [`DWIDTH-1:0] b23_data_delayed_14;
wire [`DWIDTH-1:0] b23_data_delayed_15;
wire [`DWIDTH-1:0] b23_data_delayed_16;
wire [`DWIDTH-1:0] b23_data_delayed_17;
wire [`DWIDTH-1:0] b23_data_delayed_18;
wire [`DWIDTH-1:0] b23_data_delayed_19;
wire [`DWIDTH-1:0] b23_data_delayed_20;
wire [`DWIDTH-1:0] b23_data_delayed_21;
wire [`DWIDTH-1:0] b23_data_delayed_22;
wire [`DWIDTH-1:0] b23_data_delayed_23;
wire [`DWIDTH-1:0] b24_data_delayed_1;
wire [`DWIDTH-1:0] b24_data_delayed_2;
wire [`DWIDTH-1:0] b24_data_delayed_3;
wire [`DWIDTH-1:0] b24_data_delayed_4;
wire [`DWIDTH-1:0] b24_data_delayed_5;
wire [`DWIDTH-1:0] b24_data_delayed_6;
wire [`DWIDTH-1:0] b24_data_delayed_7;
wire [`DWIDTH-1:0] b24_data_delayed_8;
wire [`DWIDTH-1:0] b24_data_delayed_9;
wire [`DWIDTH-1:0] b24_data_delayed_10;
wire [`DWIDTH-1:0] b24_data_delayed_11;
wire [`DWIDTH-1:0] b24_data_delayed_12;
wire [`DWIDTH-1:0] b24_data_delayed_13;
wire [`DWIDTH-1:0] b24_data_delayed_14;
wire [`DWIDTH-1:0] b24_data_delayed_15;
wire [`DWIDTH-1:0] b24_data_delayed_16;
wire [`DWIDTH-1:0] b24_data_delayed_17;
wire [`DWIDTH-1:0] b24_data_delayed_18;
wire [`DWIDTH-1:0] b24_data_delayed_19;
wire [`DWIDTH-1:0] b24_data_delayed_20;
wire [`DWIDTH-1:0] b24_data_delayed_21;
wire [`DWIDTH-1:0] b24_data_delayed_22;
wire [`DWIDTH-1:0] b24_data_delayed_23;
wire [`DWIDTH-1:0] b24_data_delayed_24;
wire [`DWIDTH-1:0] b25_data_delayed_1;
wire [`DWIDTH-1:0] b25_data_delayed_2;
wire [`DWIDTH-1:0] b25_data_delayed_3;
wire [`DWIDTH-1:0] b25_data_delayed_4;
wire [`DWIDTH-1:0] b25_data_delayed_5;
wire [`DWIDTH-1:0] b25_data_delayed_6;
wire [`DWIDTH-1:0] b25_data_delayed_7;
wire [`DWIDTH-1:0] b25_data_delayed_8;
wire [`DWIDTH-1:0] b25_data_delayed_9;
wire [`DWIDTH-1:0] b25_data_delayed_10;
wire [`DWIDTH-1:0] b25_data_delayed_11;
wire [`DWIDTH-1:0] b25_data_delayed_12;
wire [`DWIDTH-1:0] b25_data_delayed_13;
wire [`DWIDTH-1:0] b25_data_delayed_14;
wire [`DWIDTH-1:0] b25_data_delayed_15;
wire [`DWIDTH-1:0] b25_data_delayed_16;
wire [`DWIDTH-1:0] b25_data_delayed_17;
wire [`DWIDTH-1:0] b25_data_delayed_18;
wire [`DWIDTH-1:0] b25_data_delayed_19;
wire [`DWIDTH-1:0] b25_data_delayed_20;
wire [`DWIDTH-1:0] b25_data_delayed_21;
wire [`DWIDTH-1:0] b25_data_delayed_22;
wire [`DWIDTH-1:0] b25_data_delayed_23;
wire [`DWIDTH-1:0] b25_data_delayed_24;
wire [`DWIDTH-1:0] b25_data_delayed_25;
wire [`DWIDTH-1:0] b26_data_delayed_1;
wire [`DWIDTH-1:0] b26_data_delayed_2;
wire [`DWIDTH-1:0] b26_data_delayed_3;
wire [`DWIDTH-1:0] b26_data_delayed_4;
wire [`DWIDTH-1:0] b26_data_delayed_5;
wire [`DWIDTH-1:0] b26_data_delayed_6;
wire [`DWIDTH-1:0] b26_data_delayed_7;
wire [`DWIDTH-1:0] b26_data_delayed_8;
wire [`DWIDTH-1:0] b26_data_delayed_9;
wire [`DWIDTH-1:0] b26_data_delayed_10;
wire [`DWIDTH-1:0] b26_data_delayed_11;
wire [`DWIDTH-1:0] b26_data_delayed_12;
wire [`DWIDTH-1:0] b26_data_delayed_13;
wire [`DWIDTH-1:0] b26_data_delayed_14;
wire [`DWIDTH-1:0] b26_data_delayed_15;
wire [`DWIDTH-1:0] b26_data_delayed_16;
wire [`DWIDTH-1:0] b26_data_delayed_17;
wire [`DWIDTH-1:0] b26_data_delayed_18;
wire [`DWIDTH-1:0] b26_data_delayed_19;
wire [`DWIDTH-1:0] b26_data_delayed_20;
wire [`DWIDTH-1:0] b26_data_delayed_21;
wire [`DWIDTH-1:0] b26_data_delayed_22;
wire [`DWIDTH-1:0] b26_data_delayed_23;
wire [`DWIDTH-1:0] b26_data_delayed_24;
wire [`DWIDTH-1:0] b26_data_delayed_25;
wire [`DWIDTH-1:0] b26_data_delayed_26;
wire [`DWIDTH-1:0] b27_data_delayed_1;
wire [`DWIDTH-1:0] b27_data_delayed_2;
wire [`DWIDTH-1:0] b27_data_delayed_3;
wire [`DWIDTH-1:0] b27_data_delayed_4;
wire [`DWIDTH-1:0] b27_data_delayed_5;
wire [`DWIDTH-1:0] b27_data_delayed_6;
wire [`DWIDTH-1:0] b27_data_delayed_7;
wire [`DWIDTH-1:0] b27_data_delayed_8;
wire [`DWIDTH-1:0] b27_data_delayed_9;
wire [`DWIDTH-1:0] b27_data_delayed_10;
wire [`DWIDTH-1:0] b27_data_delayed_11;
wire [`DWIDTH-1:0] b27_data_delayed_12;
wire [`DWIDTH-1:0] b27_data_delayed_13;
wire [`DWIDTH-1:0] b27_data_delayed_14;
wire [`DWIDTH-1:0] b27_data_delayed_15;
wire [`DWIDTH-1:0] b27_data_delayed_16;
wire [`DWIDTH-1:0] b27_data_delayed_17;
wire [`DWIDTH-1:0] b27_data_delayed_18;
wire [`DWIDTH-1:0] b27_data_delayed_19;
wire [`DWIDTH-1:0] b27_data_delayed_20;
wire [`DWIDTH-1:0] b27_data_delayed_21;
wire [`DWIDTH-1:0] b27_data_delayed_22;
wire [`DWIDTH-1:0] b27_data_delayed_23;
wire [`DWIDTH-1:0] b27_data_delayed_24;
wire [`DWIDTH-1:0] b27_data_delayed_25;
wire [`DWIDTH-1:0] b27_data_delayed_26;
wire [`DWIDTH-1:0] b27_data_delayed_27;
wire [`DWIDTH-1:0] b28_data_delayed_1;
wire [`DWIDTH-1:0] b28_data_delayed_2;
wire [`DWIDTH-1:0] b28_data_delayed_3;
wire [`DWIDTH-1:0] b28_data_delayed_4;
wire [`DWIDTH-1:0] b28_data_delayed_5;
wire [`DWIDTH-1:0] b28_data_delayed_6;
wire [`DWIDTH-1:0] b28_data_delayed_7;
wire [`DWIDTH-1:0] b28_data_delayed_8;
wire [`DWIDTH-1:0] b28_data_delayed_9;
wire [`DWIDTH-1:0] b28_data_delayed_10;
wire [`DWIDTH-1:0] b28_data_delayed_11;
wire [`DWIDTH-1:0] b28_data_delayed_12;
wire [`DWIDTH-1:0] b28_data_delayed_13;
wire [`DWIDTH-1:0] b28_data_delayed_14;
wire [`DWIDTH-1:0] b28_data_delayed_15;
wire [`DWIDTH-1:0] b28_data_delayed_16;
wire [`DWIDTH-1:0] b28_data_delayed_17;
wire [`DWIDTH-1:0] b28_data_delayed_18;
wire [`DWIDTH-1:0] b28_data_delayed_19;
wire [`DWIDTH-1:0] b28_data_delayed_20;
wire [`DWIDTH-1:0] b28_data_delayed_21;
wire [`DWIDTH-1:0] b28_data_delayed_22;
wire [`DWIDTH-1:0] b28_data_delayed_23;
wire [`DWIDTH-1:0] b28_data_delayed_24;
wire [`DWIDTH-1:0] b28_data_delayed_25;
wire [`DWIDTH-1:0] b28_data_delayed_26;
wire [`DWIDTH-1:0] b28_data_delayed_27;
wire [`DWIDTH-1:0] b28_data_delayed_28;
wire [`DWIDTH-1:0] b29_data_delayed_1;
wire [`DWIDTH-1:0] b29_data_delayed_2;
wire [`DWIDTH-1:0] b29_data_delayed_3;
wire [`DWIDTH-1:0] b29_data_delayed_4;
wire [`DWIDTH-1:0] b29_data_delayed_5;
wire [`DWIDTH-1:0] b29_data_delayed_6;
wire [`DWIDTH-1:0] b29_data_delayed_7;
wire [`DWIDTH-1:0] b29_data_delayed_8;
wire [`DWIDTH-1:0] b29_data_delayed_9;
wire [`DWIDTH-1:0] b29_data_delayed_10;
wire [`DWIDTH-1:0] b29_data_delayed_11;
wire [`DWIDTH-1:0] b29_data_delayed_12;
wire [`DWIDTH-1:0] b29_data_delayed_13;
wire [`DWIDTH-1:0] b29_data_delayed_14;
wire [`DWIDTH-1:0] b29_data_delayed_15;
wire [`DWIDTH-1:0] b29_data_delayed_16;
wire [`DWIDTH-1:0] b29_data_delayed_17;
wire [`DWIDTH-1:0] b29_data_delayed_18;
wire [`DWIDTH-1:0] b29_data_delayed_19;
wire [`DWIDTH-1:0] b29_data_delayed_20;
wire [`DWIDTH-1:0] b29_data_delayed_21;
wire [`DWIDTH-1:0] b29_data_delayed_22;
wire [`DWIDTH-1:0] b29_data_delayed_23;
wire [`DWIDTH-1:0] b29_data_delayed_24;
wire [`DWIDTH-1:0] b29_data_delayed_25;
wire [`DWIDTH-1:0] b29_data_delayed_26;
wire [`DWIDTH-1:0] b29_data_delayed_27;
wire [`DWIDTH-1:0] b29_data_delayed_28;
wire [`DWIDTH-1:0] b29_data_delayed_29;
wire [`DWIDTH-1:0] b30_data_delayed_1;
wire [`DWIDTH-1:0] b30_data_delayed_2;
wire [`DWIDTH-1:0] b30_data_delayed_3;
wire [`DWIDTH-1:0] b30_data_delayed_4;
wire [`DWIDTH-1:0] b30_data_delayed_5;
wire [`DWIDTH-1:0] b30_data_delayed_6;
wire [`DWIDTH-1:0] b30_data_delayed_7;
wire [`DWIDTH-1:0] b30_data_delayed_8;
wire [`DWIDTH-1:0] b30_data_delayed_9;
wire [`DWIDTH-1:0] b30_data_delayed_10;
wire [`DWIDTH-1:0] b30_data_delayed_11;
wire [`DWIDTH-1:0] b30_data_delayed_12;
wire [`DWIDTH-1:0] b30_data_delayed_13;
wire [`DWIDTH-1:0] b30_data_delayed_14;
wire [`DWIDTH-1:0] b30_data_delayed_15;
wire [`DWIDTH-1:0] b30_data_delayed_16;
wire [`DWIDTH-1:0] b30_data_delayed_17;
wire [`DWIDTH-1:0] b30_data_delayed_18;
wire [`DWIDTH-1:0] b30_data_delayed_19;
wire [`DWIDTH-1:0] b30_data_delayed_20;
wire [`DWIDTH-1:0] b30_data_delayed_21;
wire [`DWIDTH-1:0] b30_data_delayed_22;
wire [`DWIDTH-1:0] b30_data_delayed_23;
wire [`DWIDTH-1:0] b30_data_delayed_24;
wire [`DWIDTH-1:0] b30_data_delayed_25;
wire [`DWIDTH-1:0] b30_data_delayed_26;
wire [`DWIDTH-1:0] b30_data_delayed_27;
wire [`DWIDTH-1:0] b30_data_delayed_28;
wire [`DWIDTH-1:0] b30_data_delayed_29;
wire [`DWIDTH-1:0] b30_data_delayed_30;
wire [`DWIDTH-1:0] b31_data_delayed_1;
wire [`DWIDTH-1:0] b31_data_delayed_2;
wire [`DWIDTH-1:0] b31_data_delayed_3;
wire [`DWIDTH-1:0] b31_data_delayed_4;
wire [`DWIDTH-1:0] b31_data_delayed_5;
wire [`DWIDTH-1:0] b31_data_delayed_6;
wire [`DWIDTH-1:0] b31_data_delayed_7;
wire [`DWIDTH-1:0] b31_data_delayed_8;
wire [`DWIDTH-1:0] b31_data_delayed_9;
wire [`DWIDTH-1:0] b31_data_delayed_10;
wire [`DWIDTH-1:0] b31_data_delayed_11;
wire [`DWIDTH-1:0] b31_data_delayed_12;
wire [`DWIDTH-1:0] b31_data_delayed_13;
wire [`DWIDTH-1:0] b31_data_delayed_14;
wire [`DWIDTH-1:0] b31_data_delayed_15;
wire [`DWIDTH-1:0] b31_data_delayed_16;
wire [`DWIDTH-1:0] b31_data_delayed_17;
wire [`DWIDTH-1:0] b31_data_delayed_18;
wire [`DWIDTH-1:0] b31_data_delayed_19;
wire [`DWIDTH-1:0] b31_data_delayed_20;
wire [`DWIDTH-1:0] b31_data_delayed_21;
wire [`DWIDTH-1:0] b31_data_delayed_22;
wire [`DWIDTH-1:0] b31_data_delayed_23;
wire [`DWIDTH-1:0] b31_data_delayed_24;
wire [`DWIDTH-1:0] b31_data_delayed_25;
wire [`DWIDTH-1:0] b31_data_delayed_26;
wire [`DWIDTH-1:0] b31_data_delayed_27;
wire [`DWIDTH-1:0] b31_data_delayed_28;
wire [`DWIDTH-1:0] b31_data_delayed_29;
wire [`DWIDTH-1:0] b31_data_delayed_30;
wire [`DWIDTH-1:0] b31_data_delayed_31;


//////////////////////////////////////////////////////////////////////////
// Instantiation of systolic data setup
//////////////////////////////////////////////////////////////////////////
systolic_data_setup u_systolic_data_setup(
.clk(clk),
.reset(reset),
.start_mat_mul(start_mat_mul),
.a_addr(a_addr),
.b_addr(b_addr),
.address_mat_a(address_mat_a),
.address_mat_b(address_mat_b),
.address_stride_a(address_stride_a),
.address_stride_b(address_stride_b),
.a_data(a_data),
.b_data(b_data),
.clk_cnt(clk_cnt),
.a0_data(a0_data),
.b0_data(b0_data),
.a1_data_delayed_1(a1_data_delayed_1),
.b1_data_delayed_1(b1_data_delayed_1),
.a2_data_delayed_2(a2_data_delayed_2),
.b2_data_delayed_2(b2_data_delayed_2),
.a3_data_delayed_3(a3_data_delayed_3),
.b3_data_delayed_3(b3_data_delayed_3),
.a4_data_delayed_4(a4_data_delayed_4),
.b4_data_delayed_4(b4_data_delayed_4),
.a5_data_delayed_5(a5_data_delayed_5),
.b5_data_delayed_5(b5_data_delayed_5),
.a6_data_delayed_6(a6_data_delayed_6),
.b6_data_delayed_6(b6_data_delayed_6),
.a7_data_delayed_7(a7_data_delayed_7),
.b7_data_delayed_7(b7_data_delayed_7),
.a8_data_delayed_8(a8_data_delayed_8),
.b8_data_delayed_8(b8_data_delayed_8),
.a9_data_delayed_9(a9_data_delayed_9),
.b9_data_delayed_9(b9_data_delayed_9),
.a10_data_delayed_10(a10_data_delayed_10),
.b10_data_delayed_10(b10_data_delayed_10),
.a11_data_delayed_11(a11_data_delayed_11),
.b11_data_delayed_11(b11_data_delayed_11),
.a12_data_delayed_12(a12_data_delayed_12),
.b12_data_delayed_12(b12_data_delayed_12),
.a13_data_delayed_13(a13_data_delayed_13),
.b13_data_delayed_13(b13_data_delayed_13),
.a14_data_delayed_14(a14_data_delayed_14),
.b14_data_delayed_14(b14_data_delayed_14),
.a15_data_delayed_15(a15_data_delayed_15),
.b15_data_delayed_15(b15_data_delayed_15),
.a16_data_delayed_16(a16_data_delayed_16),
.b16_data_delayed_16(b16_data_delayed_16),
.a17_data_delayed_17(a17_data_delayed_17),
.b17_data_delayed_17(b17_data_delayed_17),
.a18_data_delayed_18(a18_data_delayed_18),
.b18_data_delayed_18(b18_data_delayed_18),
.a19_data_delayed_19(a19_data_delayed_19),
.b19_data_delayed_19(b19_data_delayed_19),
.a20_data_delayed_20(a20_data_delayed_20),
.b20_data_delayed_20(b20_data_delayed_20),
.a21_data_delayed_21(a21_data_delayed_21),
.b21_data_delayed_21(b21_data_delayed_21),
.a22_data_delayed_22(a22_data_delayed_22),
.b22_data_delayed_22(b22_data_delayed_22),
.a23_data_delayed_23(a23_data_delayed_23),
.b23_data_delayed_23(b23_data_delayed_23),
.a24_data_delayed_24(a24_data_delayed_24),
.b24_data_delayed_24(b24_data_delayed_24),
.a25_data_delayed_25(a25_data_delayed_25),
.b25_data_delayed_25(b25_data_delayed_25),
.a26_data_delayed_26(a26_data_delayed_26),
.b26_data_delayed_26(b26_data_delayed_26),
.a27_data_delayed_27(a27_data_delayed_27),
.b27_data_delayed_27(b27_data_delayed_27),
.a28_data_delayed_28(a28_data_delayed_28),
.b28_data_delayed_28(b28_data_delayed_28),
.a29_data_delayed_29(a29_data_delayed_29),
.b29_data_delayed_29(b29_data_delayed_29),
.a30_data_delayed_30(a30_data_delayed_30),
.b30_data_delayed_30(b30_data_delayed_30),
.a31_data_delayed_31(a31_data_delayed_31),
.b31_data_delayed_31(b31_data_delayed_31),

.validity_mask_a_rows(validity_mask_a_rows),
.validity_mask_a_cols_b_rows(validity_mask_a_cols_b_rows),
.validity_mask_b_cols(validity_mask_b_cols),

.final_mat_mul_size(final_mat_mul_size),
  
.a_loc(a_loc),
.b_loc(b_loc)
);

//////////////////////////////////////////////////////////////////////////
// Logic to mux data_in coming from neighboring matmuls
//////////////////////////////////////////////////////////////////////////
wire [`DWIDTH-1:0] a0;
wire [`DWIDTH-1:0] a1;
wire [`DWIDTH-1:0] a2;
wire [`DWIDTH-1:0] a3;
wire [`DWIDTH-1:0] a4;
wire [`DWIDTH-1:0] a5;
wire [`DWIDTH-1:0] a6;
wire [`DWIDTH-1:0] a7;
wire [`DWIDTH-1:0] a8;
wire [`DWIDTH-1:0] a9;
wire [`DWIDTH-1:0] a10;
wire [`DWIDTH-1:0] a11;
wire [`DWIDTH-1:0] a12;
wire [`DWIDTH-1:0] a13;
wire [`DWIDTH-1:0] a14;
wire [`DWIDTH-1:0] a15;
wire [`DWIDTH-1:0] a16;
wire [`DWIDTH-1:0] a17;
wire [`DWIDTH-1:0] a18;
wire [`DWIDTH-1:0] a19;
wire [`DWIDTH-1:0] a20;
wire [`DWIDTH-1:0] a21;
wire [`DWIDTH-1:0] a22;
wire [`DWIDTH-1:0] a23;
wire [`DWIDTH-1:0] a24;
wire [`DWIDTH-1:0] a25;
wire [`DWIDTH-1:0] a26;
wire [`DWIDTH-1:0] a27;
wire [`DWIDTH-1:0] a28;
wire [`DWIDTH-1:0] a29;
wire [`DWIDTH-1:0] a30;
wire [`DWIDTH-1:0] a31;
wire [`DWIDTH-1:0] b0;
wire [`DWIDTH-1:0] b1;
wire [`DWIDTH-1:0] b2;
wire [`DWIDTH-1:0] b3;
wire [`DWIDTH-1:0] b4;
wire [`DWIDTH-1:0] b5;
wire [`DWIDTH-1:0] b6;
wire [`DWIDTH-1:0] b7;
wire [`DWIDTH-1:0] b8;
wire [`DWIDTH-1:0] b9;
wire [`DWIDTH-1:0] b10;
wire [`DWIDTH-1:0] b11;
wire [`DWIDTH-1:0] b12;
wire [`DWIDTH-1:0] b13;
wire [`DWIDTH-1:0] b14;
wire [`DWIDTH-1:0] b15;
wire [`DWIDTH-1:0] b16;
wire [`DWIDTH-1:0] b17;
wire [`DWIDTH-1:0] b18;
wire [`DWIDTH-1:0] b19;
wire [`DWIDTH-1:0] b20;
wire [`DWIDTH-1:0] b21;
wire [`DWIDTH-1:0] b22;
wire [`DWIDTH-1:0] b23;
wire [`DWIDTH-1:0] b24;
wire [`DWIDTH-1:0] b25;
wire [`DWIDTH-1:0] b26;
wire [`DWIDTH-1:0] b27;
wire [`DWIDTH-1:0] b28;
wire [`DWIDTH-1:0] b29;
wire [`DWIDTH-1:0] b30;
wire [`DWIDTH-1:0] b31;

wire [`DWIDTH-1:0] a0_data_in;
wire [`DWIDTH-1:0] a1_data_in;
wire [`DWIDTH-1:0] a2_data_in;
wire [`DWIDTH-1:0] a3_data_in;
wire [`DWIDTH-1:0] a4_data_in;
wire [`DWIDTH-1:0] a5_data_in;
wire [`DWIDTH-1:0] a6_data_in;
wire [`DWIDTH-1:0] a7_data_in;
wire [`DWIDTH-1:0] a8_data_in;
wire [`DWIDTH-1:0] a9_data_in;
wire [`DWIDTH-1:0] a10_data_in;
wire [`DWIDTH-1:0] a11_data_in;
wire [`DWIDTH-1:0] a12_data_in;
wire [`DWIDTH-1:0] a13_data_in;
wire [`DWIDTH-1:0] a14_data_in;
wire [`DWIDTH-1:0] a15_data_in;
wire [`DWIDTH-1:0] a16_data_in;
wire [`DWIDTH-1:0] a17_data_in;
wire [`DWIDTH-1:0] a18_data_in;
wire [`DWIDTH-1:0] a19_data_in;
wire [`DWIDTH-1:0] a20_data_in;
wire [`DWIDTH-1:0] a21_data_in;
wire [`DWIDTH-1:0] a22_data_in;
wire [`DWIDTH-1:0] a23_data_in;
wire [`DWIDTH-1:0] a24_data_in;
wire [`DWIDTH-1:0] a25_data_in;
wire [`DWIDTH-1:0] a26_data_in;
wire [`DWIDTH-1:0] a27_data_in;
wire [`DWIDTH-1:0] a28_data_in;
wire [`DWIDTH-1:0] a29_data_in;
wire [`DWIDTH-1:0] a30_data_in;
wire [`DWIDTH-1:0] a31_data_in;

assign a0_data_in = a_data_in[1*`DWIDTH-1:0*`DWIDTH];
assign a1_data_in = a_data_in[2*`DWIDTH-1:1*`DWIDTH];
assign a2_data_in = a_data_in[3*`DWIDTH-1:2*`DWIDTH];
assign a3_data_in = a_data_in[4*`DWIDTH-1:3*`DWIDTH];
assign a4_data_in = a_data_in[5*`DWIDTH-1:4*`DWIDTH];
assign a5_data_in = a_data_in[6*`DWIDTH-1:5*`DWIDTH];
assign a6_data_in = a_data_in[7*`DWIDTH-1:6*`DWIDTH];
assign a7_data_in = a_data_in[8*`DWIDTH-1:7*`DWIDTH];
assign a8_data_in = a_data_in[9*`DWIDTH-1:8*`DWIDTH];
assign a9_data_in = a_data_in[10*`DWIDTH-1:9*`DWIDTH];
assign a10_data_in = a_data_in[11*`DWIDTH-1:10*`DWIDTH];
assign a11_data_in = a_data_in[12*`DWIDTH-1:11*`DWIDTH];
assign a12_data_in = a_data_in[13*`DWIDTH-1:12*`DWIDTH];
assign a13_data_in = a_data_in[14*`DWIDTH-1:13*`DWIDTH];
assign a14_data_in = a_data_in[15*`DWIDTH-1:14*`DWIDTH];
assign a15_data_in = a_data_in[16*`DWIDTH-1:15*`DWIDTH];
assign a16_data_in = a_data_in[17*`DWIDTH-1:16*`DWIDTH];
assign a17_data_in = a_data_in[18*`DWIDTH-1:17*`DWIDTH];
assign a18_data_in = a_data_in[19*`DWIDTH-1:18*`DWIDTH];
assign a19_data_in = a_data_in[20*`DWIDTH-1:19*`DWIDTH];
assign a20_data_in = a_data_in[21*`DWIDTH-1:20*`DWIDTH];
assign a21_data_in = a_data_in[22*`DWIDTH-1:21*`DWIDTH];
assign a22_data_in = a_data_in[23*`DWIDTH-1:22*`DWIDTH];
assign a23_data_in = a_data_in[24*`DWIDTH-1:23*`DWIDTH];
assign a24_data_in = a_data_in[25*`DWIDTH-1:24*`DWIDTH];
assign a25_data_in = a_data_in[26*`DWIDTH-1:25*`DWIDTH];
assign a26_data_in = a_data_in[27*`DWIDTH-1:26*`DWIDTH];
assign a27_data_in = a_data_in[28*`DWIDTH-1:27*`DWIDTH];
assign a28_data_in = a_data_in[29*`DWIDTH-1:28*`DWIDTH];
assign a29_data_in = a_data_in[30*`DWIDTH-1:29*`DWIDTH];
assign a30_data_in = a_data_in[31*`DWIDTH-1:30*`DWIDTH];
assign a31_data_in = a_data_in[32*`DWIDTH-1:31*`DWIDTH];

wire [`DWIDTH-1:0] b0_data_in;
wire [`DWIDTH-1:0] b1_data_in;
wire [`DWIDTH-1:0] b2_data_in;
wire [`DWIDTH-1:0] b3_data_in;
wire [`DWIDTH-1:0] b4_data_in;
wire [`DWIDTH-1:0] b5_data_in;
wire [`DWIDTH-1:0] b6_data_in;
wire [`DWIDTH-1:0] b7_data_in;
wire [`DWIDTH-1:0] b8_data_in;
wire [`DWIDTH-1:0] b9_data_in;
wire [`DWIDTH-1:0] b10_data_in;
wire [`DWIDTH-1:0] b11_data_in;
wire [`DWIDTH-1:0] b12_data_in;
wire [`DWIDTH-1:0] b13_data_in;
wire [`DWIDTH-1:0] b14_data_in;
wire [`DWIDTH-1:0] b15_data_in;
wire [`DWIDTH-1:0] b16_data_in;
wire [`DWIDTH-1:0] b17_data_in;
wire [`DWIDTH-1:0] b18_data_in;
wire [`DWIDTH-1:0] b19_data_in;
wire [`DWIDTH-1:0] b20_data_in;
wire [`DWIDTH-1:0] b21_data_in;
wire [`DWIDTH-1:0] b22_data_in;
wire [`DWIDTH-1:0] b23_data_in;
wire [`DWIDTH-1:0] b24_data_in;
wire [`DWIDTH-1:0] b25_data_in;
wire [`DWIDTH-1:0] b26_data_in;
wire [`DWIDTH-1:0] b27_data_in;
wire [`DWIDTH-1:0] b28_data_in;
wire [`DWIDTH-1:0] b29_data_in;
wire [`DWIDTH-1:0] b30_data_in;
wire [`DWIDTH-1:0] b31_data_in;

assign b0_data_in = b_data_in[1*`DWIDTH-1:0*`DWIDTH];
assign b1_data_in = b_data_in[2*`DWIDTH-1:1*`DWIDTH];
assign b2_data_in = b_data_in[3*`DWIDTH-1:2*`DWIDTH];
assign b3_data_in = b_data_in[4*`DWIDTH-1:3*`DWIDTH];
assign b4_data_in = b_data_in[5*`DWIDTH-1:4*`DWIDTH];
assign b5_data_in = b_data_in[6*`DWIDTH-1:5*`DWIDTH];
assign b6_data_in = b_data_in[7*`DWIDTH-1:6*`DWIDTH];
assign b7_data_in = b_data_in[8*`DWIDTH-1:7*`DWIDTH];
assign b8_data_in = b_data_in[9*`DWIDTH-1:8*`DWIDTH];
assign b9_data_in = b_data_in[10*`DWIDTH-1:9*`DWIDTH];
assign b10_data_in = b_data_in[11*`DWIDTH-1:10*`DWIDTH];
assign b11_data_in = b_data_in[12*`DWIDTH-1:11*`DWIDTH];
assign b12_data_in = b_data_in[13*`DWIDTH-1:12*`DWIDTH];
assign b13_data_in = b_data_in[14*`DWIDTH-1:13*`DWIDTH];
assign b14_data_in = b_data_in[15*`DWIDTH-1:14*`DWIDTH];
assign b15_data_in = b_data_in[16*`DWIDTH-1:15*`DWIDTH];
assign b16_data_in = b_data_in[17*`DWIDTH-1:16*`DWIDTH];
assign b17_data_in = b_data_in[18*`DWIDTH-1:17*`DWIDTH];
assign b18_data_in = b_data_in[19*`DWIDTH-1:18*`DWIDTH];
assign b19_data_in = b_data_in[20*`DWIDTH-1:19*`DWIDTH];
assign b20_data_in = b_data_in[21*`DWIDTH-1:20*`DWIDTH];
assign b21_data_in = b_data_in[22*`DWIDTH-1:21*`DWIDTH];
assign b22_data_in = b_data_in[23*`DWIDTH-1:22*`DWIDTH];
assign b23_data_in = b_data_in[24*`DWIDTH-1:23*`DWIDTH];
assign b24_data_in = b_data_in[25*`DWIDTH-1:24*`DWIDTH];
assign b25_data_in = b_data_in[26*`DWIDTH-1:25*`DWIDTH];
assign b26_data_in = b_data_in[27*`DWIDTH-1:26*`DWIDTH];
assign b27_data_in = b_data_in[28*`DWIDTH-1:27*`DWIDTH];
assign b28_data_in = b_data_in[29*`DWIDTH-1:28*`DWIDTH];
assign b29_data_in = b_data_in[30*`DWIDTH-1:29*`DWIDTH];
assign b30_data_in = b_data_in[31*`DWIDTH-1:30*`DWIDTH];
assign b31_data_in = b_data_in[32*`DWIDTH-1:31*`DWIDTH];

assign a0 = (b_loc==0) ? a0_data           : a0_data_in;
assign a1 = (b_loc==0) ? a1_data_delayed_1 : a1_data_in;
assign a2 = (b_loc==0) ? a2_data_delayed_2 : a2_data_in;
assign a3 = (b_loc==0) ? a3_data_delayed_3 : a3_data_in;
assign a4 = (b_loc==0) ? a4_data_delayed_4 : a4_data_in;
assign a5 = (b_loc==0) ? a5_data_delayed_5 : a5_data_in;
assign a6 = (b_loc==0) ? a6_data_delayed_6 : a6_data_in;
assign a7 = (b_loc==0) ? a7_data_delayed_7 : a7_data_in;
assign a8 = (b_loc==0) ? a8_data_delayed_8 : a8_data_in;
assign a9 = (b_loc==0) ? a9_data_delayed_9 : a9_data_in;
assign a10 = (b_loc==0) ? a10_data_delayed_10 : a10_data_in;
assign a11 = (b_loc==0) ? a11_data_delayed_11 : a11_data_in;
assign a12 = (b_loc==0) ? a12_data_delayed_12 : a12_data_in;
assign a13 = (b_loc==0) ? a13_data_delayed_13 : a13_data_in;
assign a14 = (b_loc==0) ? a14_data_delayed_14 : a14_data_in;
assign a15 = (b_loc==0) ? a15_data_delayed_15 : a15_data_in;
assign a16 = (b_loc==0) ? a16_data_delayed_16 : a16_data_in;
assign a17 = (b_loc==0) ? a17_data_delayed_17 : a17_data_in;
assign a18 = (b_loc==0) ? a18_data_delayed_18 : a18_data_in;
assign a19 = (b_loc==0) ? a19_data_delayed_19 : a19_data_in;
assign a20 = (b_loc==0) ? a20_data_delayed_20 : a20_data_in;
assign a21 = (b_loc==0) ? a21_data_delayed_21 : a21_data_in;
assign a22 = (b_loc==0) ? a22_data_delayed_22 : a22_data_in;
assign a23 = (b_loc==0) ? a23_data_delayed_23 : a23_data_in;
assign a24 = (b_loc==0) ? a24_data_delayed_24 : a24_data_in;
assign a25 = (b_loc==0) ? a25_data_delayed_25 : a25_data_in;
assign a26 = (b_loc==0) ? a26_data_delayed_26 : a26_data_in;
assign a27 = (b_loc==0) ? a27_data_delayed_27 : a27_data_in;
assign a28 = (b_loc==0) ? a28_data_delayed_28 : a28_data_in;
assign a29 = (b_loc==0) ? a29_data_delayed_29 : a29_data_in;
assign a30 = (b_loc==0) ? a30_data_delayed_30 : a30_data_in;
assign a31 = (b_loc==0) ? a31_data_delayed_31 : a31_data_in;

assign b0 = (a_loc==0) ? b0_data           : b0_data_in;
assign b1 = (a_loc==0) ? b1_data_delayed_1 : b1_data_in;
assign b2 = (a_loc==0) ? b2_data_delayed_2 : b2_data_in;
assign b3 = (a_loc==0) ? b3_data_delayed_3 : b3_data_in;
assign b4 = (a_loc==0) ? b4_data_delayed_4 : b4_data_in;
assign b5 = (a_loc==0) ? b5_data_delayed_5 : b5_data_in;
assign b6 = (a_loc==0) ? b6_data_delayed_6 : b6_data_in;
assign b7 = (a_loc==0) ? b7_data_delayed_7 : b7_data_in;
assign b8 = (a_loc==0) ? b8_data_delayed_8 : b8_data_in;
assign b9 = (a_loc==0) ? b9_data_delayed_9 : b9_data_in;
assign b10 = (a_loc==0) ? b10_data_delayed_10 : b10_data_in;
assign b11 = (a_loc==0) ? b11_data_delayed_11 : b11_data_in;
assign b12 = (a_loc==0) ? b12_data_delayed_12 : b12_data_in;
assign b13 = (a_loc==0) ? b13_data_delayed_13 : b13_data_in;
assign b14 = (a_loc==0) ? b14_data_delayed_14 : b14_data_in;
assign b15 = (a_loc==0) ? b15_data_delayed_15 : b15_data_in;
assign b16 = (a_loc==0) ? b16_data_delayed_16 : b16_data_in;
assign b17 = (a_loc==0) ? b17_data_delayed_17 : b17_data_in;
assign b18 = (a_loc==0) ? b18_data_delayed_18 : b18_data_in;
assign b19 = (a_loc==0) ? b19_data_delayed_19 : b19_data_in;
assign b20 = (a_loc==0) ? b20_data_delayed_20 : b20_data_in;
assign b21 = (a_loc==0) ? b21_data_delayed_21 : b21_data_in;
assign b22 = (a_loc==0) ? b22_data_delayed_22 : b22_data_in;
assign b23 = (a_loc==0) ? b23_data_delayed_23 : b23_data_in;
assign b24 = (a_loc==0) ? b24_data_delayed_24 : b24_data_in;
assign b25 = (a_loc==0) ? b25_data_delayed_25 : b25_data_in;
assign b26 = (a_loc==0) ? b26_data_delayed_26 : b26_data_in;
assign b27 = (a_loc==0) ? b27_data_delayed_27 : b27_data_in;
assign b28 = (a_loc==0) ? b28_data_delayed_28 : b28_data_in;
assign b29 = (a_loc==0) ? b29_data_delayed_29 : b29_data_in;
assign b30 = (a_loc==0) ? b30_data_delayed_30 : b30_data_in;
assign b31 = (a_loc==0) ? b31_data_delayed_31 : b31_data_in;

wire [`DWIDTH-1:0] matrixC0_0;
wire [`DWIDTH-1:0] matrixC0_1;
wire [`DWIDTH-1:0] matrixC0_2;
wire [`DWIDTH-1:0] matrixC0_3;
wire [`DWIDTH-1:0] matrixC0_4;
wire [`DWIDTH-1:0] matrixC0_5;
wire [`DWIDTH-1:0] matrixC0_6;
wire [`DWIDTH-1:0] matrixC0_7;
wire [`DWIDTH-1:0] matrixC0_8;
wire [`DWIDTH-1:0] matrixC0_9;
wire [`DWIDTH-1:0] matrixC0_10;
wire [`DWIDTH-1:0] matrixC0_11;
wire [`DWIDTH-1:0] matrixC0_12;
wire [`DWIDTH-1:0] matrixC0_13;
wire [`DWIDTH-1:0] matrixC0_14;
wire [`DWIDTH-1:0] matrixC0_15;
wire [`DWIDTH-1:0] matrixC0_16;
wire [`DWIDTH-1:0] matrixC0_17;
wire [`DWIDTH-1:0] matrixC0_18;
wire [`DWIDTH-1:0] matrixC0_19;
wire [`DWIDTH-1:0] matrixC0_20;
wire [`DWIDTH-1:0] matrixC0_21;
wire [`DWIDTH-1:0] matrixC0_22;
wire [`DWIDTH-1:0] matrixC0_23;
wire [`DWIDTH-1:0] matrixC0_24;
wire [`DWIDTH-1:0] matrixC0_25;
wire [`DWIDTH-1:0] matrixC0_26;
wire [`DWIDTH-1:0] matrixC0_27;
wire [`DWIDTH-1:0] matrixC0_28;
wire [`DWIDTH-1:0] matrixC0_29;
wire [`DWIDTH-1:0] matrixC0_30;
wire [`DWIDTH-1:0] matrixC0_31;
wire [`DWIDTH-1:0] matrixC1_0;
wire [`DWIDTH-1:0] matrixC1_1;
wire [`DWIDTH-1:0] matrixC1_2;
wire [`DWIDTH-1:0] matrixC1_3;
wire [`DWIDTH-1:0] matrixC1_4;
wire [`DWIDTH-1:0] matrixC1_5;
wire [`DWIDTH-1:0] matrixC1_6;
wire [`DWIDTH-1:0] matrixC1_7;
wire [`DWIDTH-1:0] matrixC1_8;
wire [`DWIDTH-1:0] matrixC1_9;
wire [`DWIDTH-1:0] matrixC1_10;
wire [`DWIDTH-1:0] matrixC1_11;
wire [`DWIDTH-1:0] matrixC1_12;
wire [`DWIDTH-1:0] matrixC1_13;
wire [`DWIDTH-1:0] matrixC1_14;
wire [`DWIDTH-1:0] matrixC1_15;
wire [`DWIDTH-1:0] matrixC1_16;
wire [`DWIDTH-1:0] matrixC1_17;
wire [`DWIDTH-1:0] matrixC1_18;
wire [`DWIDTH-1:0] matrixC1_19;
wire [`DWIDTH-1:0] matrixC1_20;
wire [`DWIDTH-1:0] matrixC1_21;
wire [`DWIDTH-1:0] matrixC1_22;
wire [`DWIDTH-1:0] matrixC1_23;
wire [`DWIDTH-1:0] matrixC1_24;
wire [`DWIDTH-1:0] matrixC1_25;
wire [`DWIDTH-1:0] matrixC1_26;
wire [`DWIDTH-1:0] matrixC1_27;
wire [`DWIDTH-1:0] matrixC1_28;
wire [`DWIDTH-1:0] matrixC1_29;
wire [`DWIDTH-1:0] matrixC1_30;
wire [`DWIDTH-1:0] matrixC1_31;
wire [`DWIDTH-1:0] matrixC2_0;
wire [`DWIDTH-1:0] matrixC2_1;
wire [`DWIDTH-1:0] matrixC2_2;
wire [`DWIDTH-1:0] matrixC2_3;
wire [`DWIDTH-1:0] matrixC2_4;
wire [`DWIDTH-1:0] matrixC2_5;
wire [`DWIDTH-1:0] matrixC2_6;
wire [`DWIDTH-1:0] matrixC2_7;
wire [`DWIDTH-1:0] matrixC2_8;
wire [`DWIDTH-1:0] matrixC2_9;
wire [`DWIDTH-1:0] matrixC2_10;
wire [`DWIDTH-1:0] matrixC2_11;
wire [`DWIDTH-1:0] matrixC2_12;
wire [`DWIDTH-1:0] matrixC2_13;
wire [`DWIDTH-1:0] matrixC2_14;
wire [`DWIDTH-1:0] matrixC2_15;
wire [`DWIDTH-1:0] matrixC2_16;
wire [`DWIDTH-1:0] matrixC2_17;
wire [`DWIDTH-1:0] matrixC2_18;
wire [`DWIDTH-1:0] matrixC2_19;
wire [`DWIDTH-1:0] matrixC2_20;
wire [`DWIDTH-1:0] matrixC2_21;
wire [`DWIDTH-1:0] matrixC2_22;
wire [`DWIDTH-1:0] matrixC2_23;
wire [`DWIDTH-1:0] matrixC2_24;
wire [`DWIDTH-1:0] matrixC2_25;
wire [`DWIDTH-1:0] matrixC2_26;
wire [`DWIDTH-1:0] matrixC2_27;
wire [`DWIDTH-1:0] matrixC2_28;
wire [`DWIDTH-1:0] matrixC2_29;
wire [`DWIDTH-1:0] matrixC2_30;
wire [`DWIDTH-1:0] matrixC2_31;
wire [`DWIDTH-1:0] matrixC3_0;
wire [`DWIDTH-1:0] matrixC3_1;
wire [`DWIDTH-1:0] matrixC3_2;
wire [`DWIDTH-1:0] matrixC3_3;
wire [`DWIDTH-1:0] matrixC3_4;
wire [`DWIDTH-1:0] matrixC3_5;
wire [`DWIDTH-1:0] matrixC3_6;
wire [`DWIDTH-1:0] matrixC3_7;
wire [`DWIDTH-1:0] matrixC3_8;
wire [`DWIDTH-1:0] matrixC3_9;
wire [`DWIDTH-1:0] matrixC3_10;
wire [`DWIDTH-1:0] matrixC3_11;
wire [`DWIDTH-1:0] matrixC3_12;
wire [`DWIDTH-1:0] matrixC3_13;
wire [`DWIDTH-1:0] matrixC3_14;
wire [`DWIDTH-1:0] matrixC3_15;
wire [`DWIDTH-1:0] matrixC3_16;
wire [`DWIDTH-1:0] matrixC3_17;
wire [`DWIDTH-1:0] matrixC3_18;
wire [`DWIDTH-1:0] matrixC3_19;
wire [`DWIDTH-1:0] matrixC3_20;
wire [`DWIDTH-1:0] matrixC3_21;
wire [`DWIDTH-1:0] matrixC3_22;
wire [`DWIDTH-1:0] matrixC3_23;
wire [`DWIDTH-1:0] matrixC3_24;
wire [`DWIDTH-1:0] matrixC3_25;
wire [`DWIDTH-1:0] matrixC3_26;
wire [`DWIDTH-1:0] matrixC3_27;
wire [`DWIDTH-1:0] matrixC3_28;
wire [`DWIDTH-1:0] matrixC3_29;
wire [`DWIDTH-1:0] matrixC3_30;
wire [`DWIDTH-1:0] matrixC3_31;
wire [`DWIDTH-1:0] matrixC4_0;
wire [`DWIDTH-1:0] matrixC4_1;
wire [`DWIDTH-1:0] matrixC4_2;
wire [`DWIDTH-1:0] matrixC4_3;
wire [`DWIDTH-1:0] matrixC4_4;
wire [`DWIDTH-1:0] matrixC4_5;
wire [`DWIDTH-1:0] matrixC4_6;
wire [`DWIDTH-1:0] matrixC4_7;
wire [`DWIDTH-1:0] matrixC4_8;
wire [`DWIDTH-1:0] matrixC4_9;
wire [`DWIDTH-1:0] matrixC4_10;
wire [`DWIDTH-1:0] matrixC4_11;
wire [`DWIDTH-1:0] matrixC4_12;
wire [`DWIDTH-1:0] matrixC4_13;
wire [`DWIDTH-1:0] matrixC4_14;
wire [`DWIDTH-1:0] matrixC4_15;
wire [`DWIDTH-1:0] matrixC4_16;
wire [`DWIDTH-1:0] matrixC4_17;
wire [`DWIDTH-1:0] matrixC4_18;
wire [`DWIDTH-1:0] matrixC4_19;
wire [`DWIDTH-1:0] matrixC4_20;
wire [`DWIDTH-1:0] matrixC4_21;
wire [`DWIDTH-1:0] matrixC4_22;
wire [`DWIDTH-1:0] matrixC4_23;
wire [`DWIDTH-1:0] matrixC4_24;
wire [`DWIDTH-1:0] matrixC4_25;
wire [`DWIDTH-1:0] matrixC4_26;
wire [`DWIDTH-1:0] matrixC4_27;
wire [`DWIDTH-1:0] matrixC4_28;
wire [`DWIDTH-1:0] matrixC4_29;
wire [`DWIDTH-1:0] matrixC4_30;
wire [`DWIDTH-1:0] matrixC4_31;
wire [`DWIDTH-1:0] matrixC5_0;
wire [`DWIDTH-1:0] matrixC5_1;
wire [`DWIDTH-1:0] matrixC5_2;
wire [`DWIDTH-1:0] matrixC5_3;
wire [`DWIDTH-1:0] matrixC5_4;
wire [`DWIDTH-1:0] matrixC5_5;
wire [`DWIDTH-1:0] matrixC5_6;
wire [`DWIDTH-1:0] matrixC5_7;
wire [`DWIDTH-1:0] matrixC5_8;
wire [`DWIDTH-1:0] matrixC5_9;
wire [`DWIDTH-1:0] matrixC5_10;
wire [`DWIDTH-1:0] matrixC5_11;
wire [`DWIDTH-1:0] matrixC5_12;
wire [`DWIDTH-1:0] matrixC5_13;
wire [`DWIDTH-1:0] matrixC5_14;
wire [`DWIDTH-1:0] matrixC5_15;
wire [`DWIDTH-1:0] matrixC5_16;
wire [`DWIDTH-1:0] matrixC5_17;
wire [`DWIDTH-1:0] matrixC5_18;
wire [`DWIDTH-1:0] matrixC5_19;
wire [`DWIDTH-1:0] matrixC5_20;
wire [`DWIDTH-1:0] matrixC5_21;
wire [`DWIDTH-1:0] matrixC5_22;
wire [`DWIDTH-1:0] matrixC5_23;
wire [`DWIDTH-1:0] matrixC5_24;
wire [`DWIDTH-1:0] matrixC5_25;
wire [`DWIDTH-1:0] matrixC5_26;
wire [`DWIDTH-1:0] matrixC5_27;
wire [`DWIDTH-1:0] matrixC5_28;
wire [`DWIDTH-1:0] matrixC5_29;
wire [`DWIDTH-1:0] matrixC5_30;
wire [`DWIDTH-1:0] matrixC5_31;
wire [`DWIDTH-1:0] matrixC6_0;
wire [`DWIDTH-1:0] matrixC6_1;
wire [`DWIDTH-1:0] matrixC6_2;
wire [`DWIDTH-1:0] matrixC6_3;
wire [`DWIDTH-1:0] matrixC6_4;
wire [`DWIDTH-1:0] matrixC6_5;
wire [`DWIDTH-1:0] matrixC6_6;
wire [`DWIDTH-1:0] matrixC6_7;
wire [`DWIDTH-1:0] matrixC6_8;
wire [`DWIDTH-1:0] matrixC6_9;
wire [`DWIDTH-1:0] matrixC6_10;
wire [`DWIDTH-1:0] matrixC6_11;
wire [`DWIDTH-1:0] matrixC6_12;
wire [`DWIDTH-1:0] matrixC6_13;
wire [`DWIDTH-1:0] matrixC6_14;
wire [`DWIDTH-1:0] matrixC6_15;
wire [`DWIDTH-1:0] matrixC6_16;
wire [`DWIDTH-1:0] matrixC6_17;
wire [`DWIDTH-1:0] matrixC6_18;
wire [`DWIDTH-1:0] matrixC6_19;
wire [`DWIDTH-1:0] matrixC6_20;
wire [`DWIDTH-1:0] matrixC6_21;
wire [`DWIDTH-1:0] matrixC6_22;
wire [`DWIDTH-1:0] matrixC6_23;
wire [`DWIDTH-1:0] matrixC6_24;
wire [`DWIDTH-1:0] matrixC6_25;
wire [`DWIDTH-1:0] matrixC6_26;
wire [`DWIDTH-1:0] matrixC6_27;
wire [`DWIDTH-1:0] matrixC6_28;
wire [`DWIDTH-1:0] matrixC6_29;
wire [`DWIDTH-1:0] matrixC6_30;
wire [`DWIDTH-1:0] matrixC6_31;
wire [`DWIDTH-1:0] matrixC7_0;
wire [`DWIDTH-1:0] matrixC7_1;
wire [`DWIDTH-1:0] matrixC7_2;
wire [`DWIDTH-1:0] matrixC7_3;
wire [`DWIDTH-1:0] matrixC7_4;
wire [`DWIDTH-1:0] matrixC7_5;
wire [`DWIDTH-1:0] matrixC7_6;
wire [`DWIDTH-1:0] matrixC7_7;
wire [`DWIDTH-1:0] matrixC7_8;
wire [`DWIDTH-1:0] matrixC7_9;
wire [`DWIDTH-1:0] matrixC7_10;
wire [`DWIDTH-1:0] matrixC7_11;
wire [`DWIDTH-1:0] matrixC7_12;
wire [`DWIDTH-1:0] matrixC7_13;
wire [`DWIDTH-1:0] matrixC7_14;
wire [`DWIDTH-1:0] matrixC7_15;
wire [`DWIDTH-1:0] matrixC7_16;
wire [`DWIDTH-1:0] matrixC7_17;
wire [`DWIDTH-1:0] matrixC7_18;
wire [`DWIDTH-1:0] matrixC7_19;
wire [`DWIDTH-1:0] matrixC7_20;
wire [`DWIDTH-1:0] matrixC7_21;
wire [`DWIDTH-1:0] matrixC7_22;
wire [`DWIDTH-1:0] matrixC7_23;
wire [`DWIDTH-1:0] matrixC7_24;
wire [`DWIDTH-1:0] matrixC7_25;
wire [`DWIDTH-1:0] matrixC7_26;
wire [`DWIDTH-1:0] matrixC7_27;
wire [`DWIDTH-1:0] matrixC7_28;
wire [`DWIDTH-1:0] matrixC7_29;
wire [`DWIDTH-1:0] matrixC7_30;
wire [`DWIDTH-1:0] matrixC7_31;
wire [`DWIDTH-1:0] matrixC8_0;
wire [`DWIDTH-1:0] matrixC8_1;
wire [`DWIDTH-1:0] matrixC8_2;
wire [`DWIDTH-1:0] matrixC8_3;
wire [`DWIDTH-1:0] matrixC8_4;
wire [`DWIDTH-1:0] matrixC8_5;
wire [`DWIDTH-1:0] matrixC8_6;
wire [`DWIDTH-1:0] matrixC8_7;
wire [`DWIDTH-1:0] matrixC8_8;
wire [`DWIDTH-1:0] matrixC8_9;
wire [`DWIDTH-1:0] matrixC8_10;
wire [`DWIDTH-1:0] matrixC8_11;
wire [`DWIDTH-1:0] matrixC8_12;
wire [`DWIDTH-1:0] matrixC8_13;
wire [`DWIDTH-1:0] matrixC8_14;
wire [`DWIDTH-1:0] matrixC8_15;
wire [`DWIDTH-1:0] matrixC8_16;
wire [`DWIDTH-1:0] matrixC8_17;
wire [`DWIDTH-1:0] matrixC8_18;
wire [`DWIDTH-1:0] matrixC8_19;
wire [`DWIDTH-1:0] matrixC8_20;
wire [`DWIDTH-1:0] matrixC8_21;
wire [`DWIDTH-1:0] matrixC8_22;
wire [`DWIDTH-1:0] matrixC8_23;
wire [`DWIDTH-1:0] matrixC8_24;
wire [`DWIDTH-1:0] matrixC8_25;
wire [`DWIDTH-1:0] matrixC8_26;
wire [`DWIDTH-1:0] matrixC8_27;
wire [`DWIDTH-1:0] matrixC8_28;
wire [`DWIDTH-1:0] matrixC8_29;
wire [`DWIDTH-1:0] matrixC8_30;
wire [`DWIDTH-1:0] matrixC8_31;
wire [`DWIDTH-1:0] matrixC9_0;
wire [`DWIDTH-1:0] matrixC9_1;
wire [`DWIDTH-1:0] matrixC9_2;
wire [`DWIDTH-1:0] matrixC9_3;
wire [`DWIDTH-1:0] matrixC9_4;
wire [`DWIDTH-1:0] matrixC9_5;
wire [`DWIDTH-1:0] matrixC9_6;
wire [`DWIDTH-1:0] matrixC9_7;
wire [`DWIDTH-1:0] matrixC9_8;
wire [`DWIDTH-1:0] matrixC9_9;
wire [`DWIDTH-1:0] matrixC9_10;
wire [`DWIDTH-1:0] matrixC9_11;
wire [`DWIDTH-1:0] matrixC9_12;
wire [`DWIDTH-1:0] matrixC9_13;
wire [`DWIDTH-1:0] matrixC9_14;
wire [`DWIDTH-1:0] matrixC9_15;
wire [`DWIDTH-1:0] matrixC9_16;
wire [`DWIDTH-1:0] matrixC9_17;
wire [`DWIDTH-1:0] matrixC9_18;
wire [`DWIDTH-1:0] matrixC9_19;
wire [`DWIDTH-1:0] matrixC9_20;
wire [`DWIDTH-1:0] matrixC9_21;
wire [`DWIDTH-1:0] matrixC9_22;
wire [`DWIDTH-1:0] matrixC9_23;
wire [`DWIDTH-1:0] matrixC9_24;
wire [`DWIDTH-1:0] matrixC9_25;
wire [`DWIDTH-1:0] matrixC9_26;
wire [`DWIDTH-1:0] matrixC9_27;
wire [`DWIDTH-1:0] matrixC9_28;
wire [`DWIDTH-1:0] matrixC9_29;
wire [`DWIDTH-1:0] matrixC9_30;
wire [`DWIDTH-1:0] matrixC9_31;
wire [`DWIDTH-1:0] matrixC10_0;
wire [`DWIDTH-1:0] matrixC10_1;
wire [`DWIDTH-1:0] matrixC10_2;
wire [`DWIDTH-1:0] matrixC10_3;
wire [`DWIDTH-1:0] matrixC10_4;
wire [`DWIDTH-1:0] matrixC10_5;
wire [`DWIDTH-1:0] matrixC10_6;
wire [`DWIDTH-1:0] matrixC10_7;
wire [`DWIDTH-1:0] matrixC10_8;
wire [`DWIDTH-1:0] matrixC10_9;
wire [`DWIDTH-1:0] matrixC10_10;
wire [`DWIDTH-1:0] matrixC10_11;
wire [`DWIDTH-1:0] matrixC10_12;
wire [`DWIDTH-1:0] matrixC10_13;
wire [`DWIDTH-1:0] matrixC10_14;
wire [`DWIDTH-1:0] matrixC10_15;
wire [`DWIDTH-1:0] matrixC10_16;
wire [`DWIDTH-1:0] matrixC10_17;
wire [`DWIDTH-1:0] matrixC10_18;
wire [`DWIDTH-1:0] matrixC10_19;
wire [`DWIDTH-1:0] matrixC10_20;
wire [`DWIDTH-1:0] matrixC10_21;
wire [`DWIDTH-1:0] matrixC10_22;
wire [`DWIDTH-1:0] matrixC10_23;
wire [`DWIDTH-1:0] matrixC10_24;
wire [`DWIDTH-1:0] matrixC10_25;
wire [`DWIDTH-1:0] matrixC10_26;
wire [`DWIDTH-1:0] matrixC10_27;
wire [`DWIDTH-1:0] matrixC10_28;
wire [`DWIDTH-1:0] matrixC10_29;
wire [`DWIDTH-1:0] matrixC10_30;
wire [`DWIDTH-1:0] matrixC10_31;
wire [`DWIDTH-1:0] matrixC11_0;
wire [`DWIDTH-1:0] matrixC11_1;
wire [`DWIDTH-1:0] matrixC11_2;
wire [`DWIDTH-1:0] matrixC11_3;
wire [`DWIDTH-1:0] matrixC11_4;
wire [`DWIDTH-1:0] matrixC11_5;
wire [`DWIDTH-1:0] matrixC11_6;
wire [`DWIDTH-1:0] matrixC11_7;
wire [`DWIDTH-1:0] matrixC11_8;
wire [`DWIDTH-1:0] matrixC11_9;
wire [`DWIDTH-1:0] matrixC11_10;
wire [`DWIDTH-1:0] matrixC11_11;
wire [`DWIDTH-1:0] matrixC11_12;
wire [`DWIDTH-1:0] matrixC11_13;
wire [`DWIDTH-1:0] matrixC11_14;
wire [`DWIDTH-1:0] matrixC11_15;
wire [`DWIDTH-1:0] matrixC11_16;
wire [`DWIDTH-1:0] matrixC11_17;
wire [`DWIDTH-1:0] matrixC11_18;
wire [`DWIDTH-1:0] matrixC11_19;
wire [`DWIDTH-1:0] matrixC11_20;
wire [`DWIDTH-1:0] matrixC11_21;
wire [`DWIDTH-1:0] matrixC11_22;
wire [`DWIDTH-1:0] matrixC11_23;
wire [`DWIDTH-1:0] matrixC11_24;
wire [`DWIDTH-1:0] matrixC11_25;
wire [`DWIDTH-1:0] matrixC11_26;
wire [`DWIDTH-1:0] matrixC11_27;
wire [`DWIDTH-1:0] matrixC11_28;
wire [`DWIDTH-1:0] matrixC11_29;
wire [`DWIDTH-1:0] matrixC11_30;
wire [`DWIDTH-1:0] matrixC11_31;
wire [`DWIDTH-1:0] matrixC12_0;
wire [`DWIDTH-1:0] matrixC12_1;
wire [`DWIDTH-1:0] matrixC12_2;
wire [`DWIDTH-1:0] matrixC12_3;
wire [`DWIDTH-1:0] matrixC12_4;
wire [`DWIDTH-1:0] matrixC12_5;
wire [`DWIDTH-1:0] matrixC12_6;
wire [`DWIDTH-1:0] matrixC12_7;
wire [`DWIDTH-1:0] matrixC12_8;
wire [`DWIDTH-1:0] matrixC12_9;
wire [`DWIDTH-1:0] matrixC12_10;
wire [`DWIDTH-1:0] matrixC12_11;
wire [`DWIDTH-1:0] matrixC12_12;
wire [`DWIDTH-1:0] matrixC12_13;
wire [`DWIDTH-1:0] matrixC12_14;
wire [`DWIDTH-1:0] matrixC12_15;
wire [`DWIDTH-1:0] matrixC12_16;
wire [`DWIDTH-1:0] matrixC12_17;
wire [`DWIDTH-1:0] matrixC12_18;
wire [`DWIDTH-1:0] matrixC12_19;
wire [`DWIDTH-1:0] matrixC12_20;
wire [`DWIDTH-1:0] matrixC12_21;
wire [`DWIDTH-1:0] matrixC12_22;
wire [`DWIDTH-1:0] matrixC12_23;
wire [`DWIDTH-1:0] matrixC12_24;
wire [`DWIDTH-1:0] matrixC12_25;
wire [`DWIDTH-1:0] matrixC12_26;
wire [`DWIDTH-1:0] matrixC12_27;
wire [`DWIDTH-1:0] matrixC12_28;
wire [`DWIDTH-1:0] matrixC12_29;
wire [`DWIDTH-1:0] matrixC12_30;
wire [`DWIDTH-1:0] matrixC12_31;
wire [`DWIDTH-1:0] matrixC13_0;
wire [`DWIDTH-1:0] matrixC13_1;
wire [`DWIDTH-1:0] matrixC13_2;
wire [`DWIDTH-1:0] matrixC13_3;
wire [`DWIDTH-1:0] matrixC13_4;
wire [`DWIDTH-1:0] matrixC13_5;
wire [`DWIDTH-1:0] matrixC13_6;
wire [`DWIDTH-1:0] matrixC13_7;
wire [`DWIDTH-1:0] matrixC13_8;
wire [`DWIDTH-1:0] matrixC13_9;
wire [`DWIDTH-1:0] matrixC13_10;
wire [`DWIDTH-1:0] matrixC13_11;
wire [`DWIDTH-1:0] matrixC13_12;
wire [`DWIDTH-1:0] matrixC13_13;
wire [`DWIDTH-1:0] matrixC13_14;
wire [`DWIDTH-1:0] matrixC13_15;
wire [`DWIDTH-1:0] matrixC13_16;
wire [`DWIDTH-1:0] matrixC13_17;
wire [`DWIDTH-1:0] matrixC13_18;
wire [`DWIDTH-1:0] matrixC13_19;
wire [`DWIDTH-1:0] matrixC13_20;
wire [`DWIDTH-1:0] matrixC13_21;
wire [`DWIDTH-1:0] matrixC13_22;
wire [`DWIDTH-1:0] matrixC13_23;
wire [`DWIDTH-1:0] matrixC13_24;
wire [`DWIDTH-1:0] matrixC13_25;
wire [`DWIDTH-1:0] matrixC13_26;
wire [`DWIDTH-1:0] matrixC13_27;
wire [`DWIDTH-1:0] matrixC13_28;
wire [`DWIDTH-1:0] matrixC13_29;
wire [`DWIDTH-1:0] matrixC13_30;
wire [`DWIDTH-1:0] matrixC13_31;
wire [`DWIDTH-1:0] matrixC14_0;
wire [`DWIDTH-1:0] matrixC14_1;
wire [`DWIDTH-1:0] matrixC14_2;
wire [`DWIDTH-1:0] matrixC14_3;
wire [`DWIDTH-1:0] matrixC14_4;
wire [`DWIDTH-1:0] matrixC14_5;
wire [`DWIDTH-1:0] matrixC14_6;
wire [`DWIDTH-1:0] matrixC14_7;
wire [`DWIDTH-1:0] matrixC14_8;
wire [`DWIDTH-1:0] matrixC14_9;
wire [`DWIDTH-1:0] matrixC14_10;
wire [`DWIDTH-1:0] matrixC14_11;
wire [`DWIDTH-1:0] matrixC14_12;
wire [`DWIDTH-1:0] matrixC14_13;
wire [`DWIDTH-1:0] matrixC14_14;
wire [`DWIDTH-1:0] matrixC14_15;
wire [`DWIDTH-1:0] matrixC14_16;
wire [`DWIDTH-1:0] matrixC14_17;
wire [`DWIDTH-1:0] matrixC14_18;
wire [`DWIDTH-1:0] matrixC14_19;
wire [`DWIDTH-1:0] matrixC14_20;
wire [`DWIDTH-1:0] matrixC14_21;
wire [`DWIDTH-1:0] matrixC14_22;
wire [`DWIDTH-1:0] matrixC14_23;
wire [`DWIDTH-1:0] matrixC14_24;
wire [`DWIDTH-1:0] matrixC14_25;
wire [`DWIDTH-1:0] matrixC14_26;
wire [`DWIDTH-1:0] matrixC14_27;
wire [`DWIDTH-1:0] matrixC14_28;
wire [`DWIDTH-1:0] matrixC14_29;
wire [`DWIDTH-1:0] matrixC14_30;
wire [`DWIDTH-1:0] matrixC14_31;
wire [`DWIDTH-1:0] matrixC15_0;
wire [`DWIDTH-1:0] matrixC15_1;
wire [`DWIDTH-1:0] matrixC15_2;
wire [`DWIDTH-1:0] matrixC15_3;
wire [`DWIDTH-1:0] matrixC15_4;
wire [`DWIDTH-1:0] matrixC15_5;
wire [`DWIDTH-1:0] matrixC15_6;
wire [`DWIDTH-1:0] matrixC15_7;
wire [`DWIDTH-1:0] matrixC15_8;
wire [`DWIDTH-1:0] matrixC15_9;
wire [`DWIDTH-1:0] matrixC15_10;
wire [`DWIDTH-1:0] matrixC15_11;
wire [`DWIDTH-1:0] matrixC15_12;
wire [`DWIDTH-1:0] matrixC15_13;
wire [`DWIDTH-1:0] matrixC15_14;
wire [`DWIDTH-1:0] matrixC15_15;
wire [`DWIDTH-1:0] matrixC15_16;
wire [`DWIDTH-1:0] matrixC15_17;
wire [`DWIDTH-1:0] matrixC15_18;
wire [`DWIDTH-1:0] matrixC15_19;
wire [`DWIDTH-1:0] matrixC15_20;
wire [`DWIDTH-1:0] matrixC15_21;
wire [`DWIDTH-1:0] matrixC15_22;
wire [`DWIDTH-1:0] matrixC15_23;
wire [`DWIDTH-1:0] matrixC15_24;
wire [`DWIDTH-1:0] matrixC15_25;
wire [`DWIDTH-1:0] matrixC15_26;
wire [`DWIDTH-1:0] matrixC15_27;
wire [`DWIDTH-1:0] matrixC15_28;
wire [`DWIDTH-1:0] matrixC15_29;
wire [`DWIDTH-1:0] matrixC15_30;
wire [`DWIDTH-1:0] matrixC15_31;
wire [`DWIDTH-1:0] matrixC16_0;
wire [`DWIDTH-1:0] matrixC16_1;
wire [`DWIDTH-1:0] matrixC16_2;
wire [`DWIDTH-1:0] matrixC16_3;
wire [`DWIDTH-1:0] matrixC16_4;
wire [`DWIDTH-1:0] matrixC16_5;
wire [`DWIDTH-1:0] matrixC16_6;
wire [`DWIDTH-1:0] matrixC16_7;
wire [`DWIDTH-1:0] matrixC16_8;
wire [`DWIDTH-1:0] matrixC16_9;
wire [`DWIDTH-1:0] matrixC16_10;
wire [`DWIDTH-1:0] matrixC16_11;
wire [`DWIDTH-1:0] matrixC16_12;
wire [`DWIDTH-1:0] matrixC16_13;
wire [`DWIDTH-1:0] matrixC16_14;
wire [`DWIDTH-1:0] matrixC16_15;
wire [`DWIDTH-1:0] matrixC16_16;
wire [`DWIDTH-1:0] matrixC16_17;
wire [`DWIDTH-1:0] matrixC16_18;
wire [`DWIDTH-1:0] matrixC16_19;
wire [`DWIDTH-1:0] matrixC16_20;
wire [`DWIDTH-1:0] matrixC16_21;
wire [`DWIDTH-1:0] matrixC16_22;
wire [`DWIDTH-1:0] matrixC16_23;
wire [`DWIDTH-1:0] matrixC16_24;
wire [`DWIDTH-1:0] matrixC16_25;
wire [`DWIDTH-1:0] matrixC16_26;
wire [`DWIDTH-1:0] matrixC16_27;
wire [`DWIDTH-1:0] matrixC16_28;
wire [`DWIDTH-1:0] matrixC16_29;
wire [`DWIDTH-1:0] matrixC16_30;
wire [`DWIDTH-1:0] matrixC16_31;
wire [`DWIDTH-1:0] matrixC17_0;
wire [`DWIDTH-1:0] matrixC17_1;
wire [`DWIDTH-1:0] matrixC17_2;
wire [`DWIDTH-1:0] matrixC17_3;
wire [`DWIDTH-1:0] matrixC17_4;
wire [`DWIDTH-1:0] matrixC17_5;
wire [`DWIDTH-1:0] matrixC17_6;
wire [`DWIDTH-1:0] matrixC17_7;
wire [`DWIDTH-1:0] matrixC17_8;
wire [`DWIDTH-1:0] matrixC17_9;
wire [`DWIDTH-1:0] matrixC17_10;
wire [`DWIDTH-1:0] matrixC17_11;
wire [`DWIDTH-1:0] matrixC17_12;
wire [`DWIDTH-1:0] matrixC17_13;
wire [`DWIDTH-1:0] matrixC17_14;
wire [`DWIDTH-1:0] matrixC17_15;
wire [`DWIDTH-1:0] matrixC17_16;
wire [`DWIDTH-1:0] matrixC17_17;
wire [`DWIDTH-1:0] matrixC17_18;
wire [`DWIDTH-1:0] matrixC17_19;
wire [`DWIDTH-1:0] matrixC17_20;
wire [`DWIDTH-1:0] matrixC17_21;
wire [`DWIDTH-1:0] matrixC17_22;
wire [`DWIDTH-1:0] matrixC17_23;
wire [`DWIDTH-1:0] matrixC17_24;
wire [`DWIDTH-1:0] matrixC17_25;
wire [`DWIDTH-1:0] matrixC17_26;
wire [`DWIDTH-1:0] matrixC17_27;
wire [`DWIDTH-1:0] matrixC17_28;
wire [`DWIDTH-1:0] matrixC17_29;
wire [`DWIDTH-1:0] matrixC17_30;
wire [`DWIDTH-1:0] matrixC17_31;
wire [`DWIDTH-1:0] matrixC18_0;
wire [`DWIDTH-1:0] matrixC18_1;
wire [`DWIDTH-1:0] matrixC18_2;
wire [`DWIDTH-1:0] matrixC18_3;
wire [`DWIDTH-1:0] matrixC18_4;
wire [`DWIDTH-1:0] matrixC18_5;
wire [`DWIDTH-1:0] matrixC18_6;
wire [`DWIDTH-1:0] matrixC18_7;
wire [`DWIDTH-1:0] matrixC18_8;
wire [`DWIDTH-1:0] matrixC18_9;
wire [`DWIDTH-1:0] matrixC18_10;
wire [`DWIDTH-1:0] matrixC18_11;
wire [`DWIDTH-1:0] matrixC18_12;
wire [`DWIDTH-1:0] matrixC18_13;
wire [`DWIDTH-1:0] matrixC18_14;
wire [`DWIDTH-1:0] matrixC18_15;
wire [`DWIDTH-1:0] matrixC18_16;
wire [`DWIDTH-1:0] matrixC18_17;
wire [`DWIDTH-1:0] matrixC18_18;
wire [`DWIDTH-1:0] matrixC18_19;
wire [`DWIDTH-1:0] matrixC18_20;
wire [`DWIDTH-1:0] matrixC18_21;
wire [`DWIDTH-1:0] matrixC18_22;
wire [`DWIDTH-1:0] matrixC18_23;
wire [`DWIDTH-1:0] matrixC18_24;
wire [`DWIDTH-1:0] matrixC18_25;
wire [`DWIDTH-1:0] matrixC18_26;
wire [`DWIDTH-1:0] matrixC18_27;
wire [`DWIDTH-1:0] matrixC18_28;
wire [`DWIDTH-1:0] matrixC18_29;
wire [`DWIDTH-1:0] matrixC18_30;
wire [`DWIDTH-1:0] matrixC18_31;
wire [`DWIDTH-1:0] matrixC19_0;
wire [`DWIDTH-1:0] matrixC19_1;
wire [`DWIDTH-1:0] matrixC19_2;
wire [`DWIDTH-1:0] matrixC19_3;
wire [`DWIDTH-1:0] matrixC19_4;
wire [`DWIDTH-1:0] matrixC19_5;
wire [`DWIDTH-1:0] matrixC19_6;
wire [`DWIDTH-1:0] matrixC19_7;
wire [`DWIDTH-1:0] matrixC19_8;
wire [`DWIDTH-1:0] matrixC19_9;
wire [`DWIDTH-1:0] matrixC19_10;
wire [`DWIDTH-1:0] matrixC19_11;
wire [`DWIDTH-1:0] matrixC19_12;
wire [`DWIDTH-1:0] matrixC19_13;
wire [`DWIDTH-1:0] matrixC19_14;
wire [`DWIDTH-1:0] matrixC19_15;
wire [`DWIDTH-1:0] matrixC19_16;
wire [`DWIDTH-1:0] matrixC19_17;
wire [`DWIDTH-1:0] matrixC19_18;
wire [`DWIDTH-1:0] matrixC19_19;
wire [`DWIDTH-1:0] matrixC19_20;
wire [`DWIDTH-1:0] matrixC19_21;
wire [`DWIDTH-1:0] matrixC19_22;
wire [`DWIDTH-1:0] matrixC19_23;
wire [`DWIDTH-1:0] matrixC19_24;
wire [`DWIDTH-1:0] matrixC19_25;
wire [`DWIDTH-1:0] matrixC19_26;
wire [`DWIDTH-1:0] matrixC19_27;
wire [`DWIDTH-1:0] matrixC19_28;
wire [`DWIDTH-1:0] matrixC19_29;
wire [`DWIDTH-1:0] matrixC19_30;
wire [`DWIDTH-1:0] matrixC19_31;
wire [`DWIDTH-1:0] matrixC20_0;
wire [`DWIDTH-1:0] matrixC20_1;
wire [`DWIDTH-1:0] matrixC20_2;
wire [`DWIDTH-1:0] matrixC20_3;
wire [`DWIDTH-1:0] matrixC20_4;
wire [`DWIDTH-1:0] matrixC20_5;
wire [`DWIDTH-1:0] matrixC20_6;
wire [`DWIDTH-1:0] matrixC20_7;
wire [`DWIDTH-1:0] matrixC20_8;
wire [`DWIDTH-1:0] matrixC20_9;
wire [`DWIDTH-1:0] matrixC20_10;
wire [`DWIDTH-1:0] matrixC20_11;
wire [`DWIDTH-1:0] matrixC20_12;
wire [`DWIDTH-1:0] matrixC20_13;
wire [`DWIDTH-1:0] matrixC20_14;
wire [`DWIDTH-1:0] matrixC20_15;
wire [`DWIDTH-1:0] matrixC20_16;
wire [`DWIDTH-1:0] matrixC20_17;
wire [`DWIDTH-1:0] matrixC20_18;
wire [`DWIDTH-1:0] matrixC20_19;
wire [`DWIDTH-1:0] matrixC20_20;
wire [`DWIDTH-1:0] matrixC20_21;
wire [`DWIDTH-1:0] matrixC20_22;
wire [`DWIDTH-1:0] matrixC20_23;
wire [`DWIDTH-1:0] matrixC20_24;
wire [`DWIDTH-1:0] matrixC20_25;
wire [`DWIDTH-1:0] matrixC20_26;
wire [`DWIDTH-1:0] matrixC20_27;
wire [`DWIDTH-1:0] matrixC20_28;
wire [`DWIDTH-1:0] matrixC20_29;
wire [`DWIDTH-1:0] matrixC20_30;
wire [`DWIDTH-1:0] matrixC20_31;
wire [`DWIDTH-1:0] matrixC21_0;
wire [`DWIDTH-1:0] matrixC21_1;
wire [`DWIDTH-1:0] matrixC21_2;
wire [`DWIDTH-1:0] matrixC21_3;
wire [`DWIDTH-1:0] matrixC21_4;
wire [`DWIDTH-1:0] matrixC21_5;
wire [`DWIDTH-1:0] matrixC21_6;
wire [`DWIDTH-1:0] matrixC21_7;
wire [`DWIDTH-1:0] matrixC21_8;
wire [`DWIDTH-1:0] matrixC21_9;
wire [`DWIDTH-1:0] matrixC21_10;
wire [`DWIDTH-1:0] matrixC21_11;
wire [`DWIDTH-1:0] matrixC21_12;
wire [`DWIDTH-1:0] matrixC21_13;
wire [`DWIDTH-1:0] matrixC21_14;
wire [`DWIDTH-1:0] matrixC21_15;
wire [`DWIDTH-1:0] matrixC21_16;
wire [`DWIDTH-1:0] matrixC21_17;
wire [`DWIDTH-1:0] matrixC21_18;
wire [`DWIDTH-1:0] matrixC21_19;
wire [`DWIDTH-1:0] matrixC21_20;
wire [`DWIDTH-1:0] matrixC21_21;
wire [`DWIDTH-1:0] matrixC21_22;
wire [`DWIDTH-1:0] matrixC21_23;
wire [`DWIDTH-1:0] matrixC21_24;
wire [`DWIDTH-1:0] matrixC21_25;
wire [`DWIDTH-1:0] matrixC21_26;
wire [`DWIDTH-1:0] matrixC21_27;
wire [`DWIDTH-1:0] matrixC21_28;
wire [`DWIDTH-1:0] matrixC21_29;
wire [`DWIDTH-1:0] matrixC21_30;
wire [`DWIDTH-1:0] matrixC21_31;
wire [`DWIDTH-1:0] matrixC22_0;
wire [`DWIDTH-1:0] matrixC22_1;
wire [`DWIDTH-1:0] matrixC22_2;
wire [`DWIDTH-1:0] matrixC22_3;
wire [`DWIDTH-1:0] matrixC22_4;
wire [`DWIDTH-1:0] matrixC22_5;
wire [`DWIDTH-1:0] matrixC22_6;
wire [`DWIDTH-1:0] matrixC22_7;
wire [`DWIDTH-1:0] matrixC22_8;
wire [`DWIDTH-1:0] matrixC22_9;
wire [`DWIDTH-1:0] matrixC22_10;
wire [`DWIDTH-1:0] matrixC22_11;
wire [`DWIDTH-1:0] matrixC22_12;
wire [`DWIDTH-1:0] matrixC22_13;
wire [`DWIDTH-1:0] matrixC22_14;
wire [`DWIDTH-1:0] matrixC22_15;
wire [`DWIDTH-1:0] matrixC22_16;
wire [`DWIDTH-1:0] matrixC22_17;
wire [`DWIDTH-1:0] matrixC22_18;
wire [`DWIDTH-1:0] matrixC22_19;
wire [`DWIDTH-1:0] matrixC22_20;
wire [`DWIDTH-1:0] matrixC22_21;
wire [`DWIDTH-1:0] matrixC22_22;
wire [`DWIDTH-1:0] matrixC22_23;
wire [`DWIDTH-1:0] matrixC22_24;
wire [`DWIDTH-1:0] matrixC22_25;
wire [`DWIDTH-1:0] matrixC22_26;
wire [`DWIDTH-1:0] matrixC22_27;
wire [`DWIDTH-1:0] matrixC22_28;
wire [`DWIDTH-1:0] matrixC22_29;
wire [`DWIDTH-1:0] matrixC22_30;
wire [`DWIDTH-1:0] matrixC22_31;
wire [`DWIDTH-1:0] matrixC23_0;
wire [`DWIDTH-1:0] matrixC23_1;
wire [`DWIDTH-1:0] matrixC23_2;
wire [`DWIDTH-1:0] matrixC23_3;
wire [`DWIDTH-1:0] matrixC23_4;
wire [`DWIDTH-1:0] matrixC23_5;
wire [`DWIDTH-1:0] matrixC23_6;
wire [`DWIDTH-1:0] matrixC23_7;
wire [`DWIDTH-1:0] matrixC23_8;
wire [`DWIDTH-1:0] matrixC23_9;
wire [`DWIDTH-1:0] matrixC23_10;
wire [`DWIDTH-1:0] matrixC23_11;
wire [`DWIDTH-1:0] matrixC23_12;
wire [`DWIDTH-1:0] matrixC23_13;
wire [`DWIDTH-1:0] matrixC23_14;
wire [`DWIDTH-1:0] matrixC23_15;
wire [`DWIDTH-1:0] matrixC23_16;
wire [`DWIDTH-1:0] matrixC23_17;
wire [`DWIDTH-1:0] matrixC23_18;
wire [`DWIDTH-1:0] matrixC23_19;
wire [`DWIDTH-1:0] matrixC23_20;
wire [`DWIDTH-1:0] matrixC23_21;
wire [`DWIDTH-1:0] matrixC23_22;
wire [`DWIDTH-1:0] matrixC23_23;
wire [`DWIDTH-1:0] matrixC23_24;
wire [`DWIDTH-1:0] matrixC23_25;
wire [`DWIDTH-1:0] matrixC23_26;
wire [`DWIDTH-1:0] matrixC23_27;
wire [`DWIDTH-1:0] matrixC23_28;
wire [`DWIDTH-1:0] matrixC23_29;
wire [`DWIDTH-1:0] matrixC23_30;
wire [`DWIDTH-1:0] matrixC23_31;
wire [`DWIDTH-1:0] matrixC24_0;
wire [`DWIDTH-1:0] matrixC24_1;
wire [`DWIDTH-1:0] matrixC24_2;
wire [`DWIDTH-1:0] matrixC24_3;
wire [`DWIDTH-1:0] matrixC24_4;
wire [`DWIDTH-1:0] matrixC24_5;
wire [`DWIDTH-1:0] matrixC24_6;
wire [`DWIDTH-1:0] matrixC24_7;
wire [`DWIDTH-1:0] matrixC24_8;
wire [`DWIDTH-1:0] matrixC24_9;
wire [`DWIDTH-1:0] matrixC24_10;
wire [`DWIDTH-1:0] matrixC24_11;
wire [`DWIDTH-1:0] matrixC24_12;
wire [`DWIDTH-1:0] matrixC24_13;
wire [`DWIDTH-1:0] matrixC24_14;
wire [`DWIDTH-1:0] matrixC24_15;
wire [`DWIDTH-1:0] matrixC24_16;
wire [`DWIDTH-1:0] matrixC24_17;
wire [`DWIDTH-1:0] matrixC24_18;
wire [`DWIDTH-1:0] matrixC24_19;
wire [`DWIDTH-1:0] matrixC24_20;
wire [`DWIDTH-1:0] matrixC24_21;
wire [`DWIDTH-1:0] matrixC24_22;
wire [`DWIDTH-1:0] matrixC24_23;
wire [`DWIDTH-1:0] matrixC24_24;
wire [`DWIDTH-1:0] matrixC24_25;
wire [`DWIDTH-1:0] matrixC24_26;
wire [`DWIDTH-1:0] matrixC24_27;
wire [`DWIDTH-1:0] matrixC24_28;
wire [`DWIDTH-1:0] matrixC24_29;
wire [`DWIDTH-1:0] matrixC24_30;
wire [`DWIDTH-1:0] matrixC24_31;
wire [`DWIDTH-1:0] matrixC25_0;
wire [`DWIDTH-1:0] matrixC25_1;
wire [`DWIDTH-1:0] matrixC25_2;
wire [`DWIDTH-1:0] matrixC25_3;
wire [`DWIDTH-1:0] matrixC25_4;
wire [`DWIDTH-1:0] matrixC25_5;
wire [`DWIDTH-1:0] matrixC25_6;
wire [`DWIDTH-1:0] matrixC25_7;
wire [`DWIDTH-1:0] matrixC25_8;
wire [`DWIDTH-1:0] matrixC25_9;
wire [`DWIDTH-1:0] matrixC25_10;
wire [`DWIDTH-1:0] matrixC25_11;
wire [`DWIDTH-1:0] matrixC25_12;
wire [`DWIDTH-1:0] matrixC25_13;
wire [`DWIDTH-1:0] matrixC25_14;
wire [`DWIDTH-1:0] matrixC25_15;
wire [`DWIDTH-1:0] matrixC25_16;
wire [`DWIDTH-1:0] matrixC25_17;
wire [`DWIDTH-1:0] matrixC25_18;
wire [`DWIDTH-1:0] matrixC25_19;
wire [`DWIDTH-1:0] matrixC25_20;
wire [`DWIDTH-1:0] matrixC25_21;
wire [`DWIDTH-1:0] matrixC25_22;
wire [`DWIDTH-1:0] matrixC25_23;
wire [`DWIDTH-1:0] matrixC25_24;
wire [`DWIDTH-1:0] matrixC25_25;
wire [`DWIDTH-1:0] matrixC25_26;
wire [`DWIDTH-1:0] matrixC25_27;
wire [`DWIDTH-1:0] matrixC25_28;
wire [`DWIDTH-1:0] matrixC25_29;
wire [`DWIDTH-1:0] matrixC25_30;
wire [`DWIDTH-1:0] matrixC25_31;
wire [`DWIDTH-1:0] matrixC26_0;
wire [`DWIDTH-1:0] matrixC26_1;
wire [`DWIDTH-1:0] matrixC26_2;
wire [`DWIDTH-1:0] matrixC26_3;
wire [`DWIDTH-1:0] matrixC26_4;
wire [`DWIDTH-1:0] matrixC26_5;
wire [`DWIDTH-1:0] matrixC26_6;
wire [`DWIDTH-1:0] matrixC26_7;
wire [`DWIDTH-1:0] matrixC26_8;
wire [`DWIDTH-1:0] matrixC26_9;
wire [`DWIDTH-1:0] matrixC26_10;
wire [`DWIDTH-1:0] matrixC26_11;
wire [`DWIDTH-1:0] matrixC26_12;
wire [`DWIDTH-1:0] matrixC26_13;
wire [`DWIDTH-1:0] matrixC26_14;
wire [`DWIDTH-1:0] matrixC26_15;
wire [`DWIDTH-1:0] matrixC26_16;
wire [`DWIDTH-1:0] matrixC26_17;
wire [`DWIDTH-1:0] matrixC26_18;
wire [`DWIDTH-1:0] matrixC26_19;
wire [`DWIDTH-1:0] matrixC26_20;
wire [`DWIDTH-1:0] matrixC26_21;
wire [`DWIDTH-1:0] matrixC26_22;
wire [`DWIDTH-1:0] matrixC26_23;
wire [`DWIDTH-1:0] matrixC26_24;
wire [`DWIDTH-1:0] matrixC26_25;
wire [`DWIDTH-1:0] matrixC26_26;
wire [`DWIDTH-1:0] matrixC26_27;
wire [`DWIDTH-1:0] matrixC26_28;
wire [`DWIDTH-1:0] matrixC26_29;
wire [`DWIDTH-1:0] matrixC26_30;
wire [`DWIDTH-1:0] matrixC26_31;
wire [`DWIDTH-1:0] matrixC27_0;
wire [`DWIDTH-1:0] matrixC27_1;
wire [`DWIDTH-1:0] matrixC27_2;
wire [`DWIDTH-1:0] matrixC27_3;
wire [`DWIDTH-1:0] matrixC27_4;
wire [`DWIDTH-1:0] matrixC27_5;
wire [`DWIDTH-1:0] matrixC27_6;
wire [`DWIDTH-1:0] matrixC27_7;
wire [`DWIDTH-1:0] matrixC27_8;
wire [`DWIDTH-1:0] matrixC27_9;
wire [`DWIDTH-1:0] matrixC27_10;
wire [`DWIDTH-1:0] matrixC27_11;
wire [`DWIDTH-1:0] matrixC27_12;
wire [`DWIDTH-1:0] matrixC27_13;
wire [`DWIDTH-1:0] matrixC27_14;
wire [`DWIDTH-1:0] matrixC27_15;
wire [`DWIDTH-1:0] matrixC27_16;
wire [`DWIDTH-1:0] matrixC27_17;
wire [`DWIDTH-1:0] matrixC27_18;
wire [`DWIDTH-1:0] matrixC27_19;
wire [`DWIDTH-1:0] matrixC27_20;
wire [`DWIDTH-1:0] matrixC27_21;
wire [`DWIDTH-1:0] matrixC27_22;
wire [`DWIDTH-1:0] matrixC27_23;
wire [`DWIDTH-1:0] matrixC27_24;
wire [`DWIDTH-1:0] matrixC27_25;
wire [`DWIDTH-1:0] matrixC27_26;
wire [`DWIDTH-1:0] matrixC27_27;
wire [`DWIDTH-1:0] matrixC27_28;
wire [`DWIDTH-1:0] matrixC27_29;
wire [`DWIDTH-1:0] matrixC27_30;
wire [`DWIDTH-1:0] matrixC27_31;
wire [`DWIDTH-1:0] matrixC28_0;
wire [`DWIDTH-1:0] matrixC28_1;
wire [`DWIDTH-1:0] matrixC28_2;
wire [`DWIDTH-1:0] matrixC28_3;
wire [`DWIDTH-1:0] matrixC28_4;
wire [`DWIDTH-1:0] matrixC28_5;
wire [`DWIDTH-1:0] matrixC28_6;
wire [`DWIDTH-1:0] matrixC28_7;
wire [`DWIDTH-1:0] matrixC28_8;
wire [`DWIDTH-1:0] matrixC28_9;
wire [`DWIDTH-1:0] matrixC28_10;
wire [`DWIDTH-1:0] matrixC28_11;
wire [`DWIDTH-1:0] matrixC28_12;
wire [`DWIDTH-1:0] matrixC28_13;
wire [`DWIDTH-1:0] matrixC28_14;
wire [`DWIDTH-1:0] matrixC28_15;
wire [`DWIDTH-1:0] matrixC28_16;
wire [`DWIDTH-1:0] matrixC28_17;
wire [`DWIDTH-1:0] matrixC28_18;
wire [`DWIDTH-1:0] matrixC28_19;
wire [`DWIDTH-1:0] matrixC28_20;
wire [`DWIDTH-1:0] matrixC28_21;
wire [`DWIDTH-1:0] matrixC28_22;
wire [`DWIDTH-1:0] matrixC28_23;
wire [`DWIDTH-1:0] matrixC28_24;
wire [`DWIDTH-1:0] matrixC28_25;
wire [`DWIDTH-1:0] matrixC28_26;
wire [`DWIDTH-1:0] matrixC28_27;
wire [`DWIDTH-1:0] matrixC28_28;
wire [`DWIDTH-1:0] matrixC28_29;
wire [`DWIDTH-1:0] matrixC28_30;
wire [`DWIDTH-1:0] matrixC28_31;
wire [`DWIDTH-1:0] matrixC29_0;
wire [`DWIDTH-1:0] matrixC29_1;
wire [`DWIDTH-1:0] matrixC29_2;
wire [`DWIDTH-1:0] matrixC29_3;
wire [`DWIDTH-1:0] matrixC29_4;
wire [`DWIDTH-1:0] matrixC29_5;
wire [`DWIDTH-1:0] matrixC29_6;
wire [`DWIDTH-1:0] matrixC29_7;
wire [`DWIDTH-1:0] matrixC29_8;
wire [`DWIDTH-1:0] matrixC29_9;
wire [`DWIDTH-1:0] matrixC29_10;
wire [`DWIDTH-1:0] matrixC29_11;
wire [`DWIDTH-1:0] matrixC29_12;
wire [`DWIDTH-1:0] matrixC29_13;
wire [`DWIDTH-1:0] matrixC29_14;
wire [`DWIDTH-1:0] matrixC29_15;
wire [`DWIDTH-1:0] matrixC29_16;
wire [`DWIDTH-1:0] matrixC29_17;
wire [`DWIDTH-1:0] matrixC29_18;
wire [`DWIDTH-1:0] matrixC29_19;
wire [`DWIDTH-1:0] matrixC29_20;
wire [`DWIDTH-1:0] matrixC29_21;
wire [`DWIDTH-1:0] matrixC29_22;
wire [`DWIDTH-1:0] matrixC29_23;
wire [`DWIDTH-1:0] matrixC29_24;
wire [`DWIDTH-1:0] matrixC29_25;
wire [`DWIDTH-1:0] matrixC29_26;
wire [`DWIDTH-1:0] matrixC29_27;
wire [`DWIDTH-1:0] matrixC29_28;
wire [`DWIDTH-1:0] matrixC29_29;
wire [`DWIDTH-1:0] matrixC29_30;
wire [`DWIDTH-1:0] matrixC29_31;
wire [`DWIDTH-1:0] matrixC30_0;
wire [`DWIDTH-1:0] matrixC30_1;
wire [`DWIDTH-1:0] matrixC30_2;
wire [`DWIDTH-1:0] matrixC30_3;
wire [`DWIDTH-1:0] matrixC30_4;
wire [`DWIDTH-1:0] matrixC30_5;
wire [`DWIDTH-1:0] matrixC30_6;
wire [`DWIDTH-1:0] matrixC30_7;
wire [`DWIDTH-1:0] matrixC30_8;
wire [`DWIDTH-1:0] matrixC30_9;
wire [`DWIDTH-1:0] matrixC30_10;
wire [`DWIDTH-1:0] matrixC30_11;
wire [`DWIDTH-1:0] matrixC30_12;
wire [`DWIDTH-1:0] matrixC30_13;
wire [`DWIDTH-1:0] matrixC30_14;
wire [`DWIDTH-1:0] matrixC30_15;
wire [`DWIDTH-1:0] matrixC30_16;
wire [`DWIDTH-1:0] matrixC30_17;
wire [`DWIDTH-1:0] matrixC30_18;
wire [`DWIDTH-1:0] matrixC30_19;
wire [`DWIDTH-1:0] matrixC30_20;
wire [`DWIDTH-1:0] matrixC30_21;
wire [`DWIDTH-1:0] matrixC30_22;
wire [`DWIDTH-1:0] matrixC30_23;
wire [`DWIDTH-1:0] matrixC30_24;
wire [`DWIDTH-1:0] matrixC30_25;
wire [`DWIDTH-1:0] matrixC30_26;
wire [`DWIDTH-1:0] matrixC30_27;
wire [`DWIDTH-1:0] matrixC30_28;
wire [`DWIDTH-1:0] matrixC30_29;
wire [`DWIDTH-1:0] matrixC30_30;
wire [`DWIDTH-1:0] matrixC30_31;
wire [`DWIDTH-1:0] matrixC31_0;
wire [`DWIDTH-1:0] matrixC31_1;
wire [`DWIDTH-1:0] matrixC31_2;
wire [`DWIDTH-1:0] matrixC31_3;
wire [`DWIDTH-1:0] matrixC31_4;
wire [`DWIDTH-1:0] matrixC31_5;
wire [`DWIDTH-1:0] matrixC31_6;
wire [`DWIDTH-1:0] matrixC31_7;
wire [`DWIDTH-1:0] matrixC31_8;
wire [`DWIDTH-1:0] matrixC31_9;
wire [`DWIDTH-1:0] matrixC31_10;
wire [`DWIDTH-1:0] matrixC31_11;
wire [`DWIDTH-1:0] matrixC31_12;
wire [`DWIDTH-1:0] matrixC31_13;
wire [`DWIDTH-1:0] matrixC31_14;
wire [`DWIDTH-1:0] matrixC31_15;
wire [`DWIDTH-1:0] matrixC31_16;
wire [`DWIDTH-1:0] matrixC31_17;
wire [`DWIDTH-1:0] matrixC31_18;
wire [`DWIDTH-1:0] matrixC31_19;
wire [`DWIDTH-1:0] matrixC31_20;
wire [`DWIDTH-1:0] matrixC31_21;
wire [`DWIDTH-1:0] matrixC31_22;
wire [`DWIDTH-1:0] matrixC31_23;
wire [`DWIDTH-1:0] matrixC31_24;
wire [`DWIDTH-1:0] matrixC31_25;
wire [`DWIDTH-1:0] matrixC31_26;
wire [`DWIDTH-1:0] matrixC31_27;
wire [`DWIDTH-1:0] matrixC31_28;
wire [`DWIDTH-1:0] matrixC31_29;
wire [`DWIDTH-1:0] matrixC31_30;
wire [`DWIDTH-1:0] matrixC31_31;


//////////////////////////////////////////////////////////////////////////
// Instantiation of the output logic
//////////////////////////////////////////////////////////////////////////
output_logic u_output_logic(
.start_mat_mul(start_mat_mul),
.done_mat_mul(done_mat_mul),
.address_mat_c(address_mat_c),
.address_stride_c(address_stride_c),
.c_data_out(c_data_out),
.c_data_in(c_data_in),
.c_addr(c_addr),
.c_data_available(c_data_available),
.clk_cnt(clk_cnt),
.row_latch_en(row_latch_en),

.final_mat_mul_size(final_mat_mul_size),
  .matrixC0_0(matrixC0_0),
.matrixC0_1(matrixC0_1),
.matrixC0_2(matrixC0_2),
.matrixC0_3(matrixC0_3),
.matrixC0_4(matrixC0_4),
.matrixC0_5(matrixC0_5),
.matrixC0_6(matrixC0_6),
.matrixC0_7(matrixC0_7),
.matrixC0_8(matrixC0_8),
.matrixC0_9(matrixC0_9),
.matrixC0_10(matrixC0_10),
.matrixC0_11(matrixC0_11),
.matrixC0_12(matrixC0_12),
.matrixC0_13(matrixC0_13),
.matrixC0_14(matrixC0_14),
.matrixC0_15(matrixC0_15),
.matrixC0_16(matrixC0_16),
.matrixC0_17(matrixC0_17),
.matrixC0_18(matrixC0_18),
.matrixC0_19(matrixC0_19),
.matrixC0_20(matrixC0_20),
.matrixC0_21(matrixC0_21),
.matrixC0_22(matrixC0_22),
.matrixC0_23(matrixC0_23),
.matrixC0_24(matrixC0_24),
.matrixC0_25(matrixC0_25),
.matrixC0_26(matrixC0_26),
.matrixC0_27(matrixC0_27),
.matrixC0_28(matrixC0_28),
.matrixC0_29(matrixC0_29),
.matrixC0_30(matrixC0_30),
.matrixC0_31(matrixC0_31),
.matrixC1_0(matrixC1_0),
.matrixC1_1(matrixC1_1),
.matrixC1_2(matrixC1_2),
.matrixC1_3(matrixC1_3),
.matrixC1_4(matrixC1_4),
.matrixC1_5(matrixC1_5),
.matrixC1_6(matrixC1_6),
.matrixC1_7(matrixC1_7),
.matrixC1_8(matrixC1_8),
.matrixC1_9(matrixC1_9),
.matrixC1_10(matrixC1_10),
.matrixC1_11(matrixC1_11),
.matrixC1_12(matrixC1_12),
.matrixC1_13(matrixC1_13),
.matrixC1_14(matrixC1_14),
.matrixC1_15(matrixC1_15),
.matrixC1_16(matrixC1_16),
.matrixC1_17(matrixC1_17),
.matrixC1_18(matrixC1_18),
.matrixC1_19(matrixC1_19),
.matrixC1_20(matrixC1_20),
.matrixC1_21(matrixC1_21),
.matrixC1_22(matrixC1_22),
.matrixC1_23(matrixC1_23),
.matrixC1_24(matrixC1_24),
.matrixC1_25(matrixC1_25),
.matrixC1_26(matrixC1_26),
.matrixC1_27(matrixC1_27),
.matrixC1_28(matrixC1_28),
.matrixC1_29(matrixC1_29),
.matrixC1_30(matrixC1_30),
.matrixC1_31(matrixC1_31),
.matrixC2_0(matrixC2_0),
.matrixC2_1(matrixC2_1),
.matrixC2_2(matrixC2_2),
.matrixC2_3(matrixC2_3),
.matrixC2_4(matrixC2_4),
.matrixC2_5(matrixC2_5),
.matrixC2_6(matrixC2_6),
.matrixC2_7(matrixC2_7),
.matrixC2_8(matrixC2_8),
.matrixC2_9(matrixC2_9),
.matrixC2_10(matrixC2_10),
.matrixC2_11(matrixC2_11),
.matrixC2_12(matrixC2_12),
.matrixC2_13(matrixC2_13),
.matrixC2_14(matrixC2_14),
.matrixC2_15(matrixC2_15),
.matrixC2_16(matrixC2_16),
.matrixC2_17(matrixC2_17),
.matrixC2_18(matrixC2_18),
.matrixC2_19(matrixC2_19),
.matrixC2_20(matrixC2_20),
.matrixC2_21(matrixC2_21),
.matrixC2_22(matrixC2_22),
.matrixC2_23(matrixC2_23),
.matrixC2_24(matrixC2_24),
.matrixC2_25(matrixC2_25),
.matrixC2_26(matrixC2_26),
.matrixC2_27(matrixC2_27),
.matrixC2_28(matrixC2_28),
.matrixC2_29(matrixC2_29),
.matrixC2_30(matrixC2_30),
.matrixC2_31(matrixC2_31),
.matrixC3_0(matrixC3_0),
.matrixC3_1(matrixC3_1),
.matrixC3_2(matrixC3_2),
.matrixC3_3(matrixC3_3),
.matrixC3_4(matrixC3_4),
.matrixC3_5(matrixC3_5),
.matrixC3_6(matrixC3_6),
.matrixC3_7(matrixC3_7),
.matrixC3_8(matrixC3_8),
.matrixC3_9(matrixC3_9),
.matrixC3_10(matrixC3_10),
.matrixC3_11(matrixC3_11),
.matrixC3_12(matrixC3_12),
.matrixC3_13(matrixC3_13),
.matrixC3_14(matrixC3_14),
.matrixC3_15(matrixC3_15),
.matrixC3_16(matrixC3_16),
.matrixC3_17(matrixC3_17),
.matrixC3_18(matrixC3_18),
.matrixC3_19(matrixC3_19),
.matrixC3_20(matrixC3_20),
.matrixC3_21(matrixC3_21),
.matrixC3_22(matrixC3_22),
.matrixC3_23(matrixC3_23),
.matrixC3_24(matrixC3_24),
.matrixC3_25(matrixC3_25),
.matrixC3_26(matrixC3_26),
.matrixC3_27(matrixC3_27),
.matrixC3_28(matrixC3_28),
.matrixC3_29(matrixC3_29),
.matrixC3_30(matrixC3_30),
.matrixC3_31(matrixC3_31),
.matrixC4_0(matrixC4_0),
.matrixC4_1(matrixC4_1),
.matrixC4_2(matrixC4_2),
.matrixC4_3(matrixC4_3),
.matrixC4_4(matrixC4_4),
.matrixC4_5(matrixC4_5),
.matrixC4_6(matrixC4_6),
.matrixC4_7(matrixC4_7),
.matrixC4_8(matrixC4_8),
.matrixC4_9(matrixC4_9),
.matrixC4_10(matrixC4_10),
.matrixC4_11(matrixC4_11),
.matrixC4_12(matrixC4_12),
.matrixC4_13(matrixC4_13),
.matrixC4_14(matrixC4_14),
.matrixC4_15(matrixC4_15),
.matrixC4_16(matrixC4_16),
.matrixC4_17(matrixC4_17),
.matrixC4_18(matrixC4_18),
.matrixC4_19(matrixC4_19),
.matrixC4_20(matrixC4_20),
.matrixC4_21(matrixC4_21),
.matrixC4_22(matrixC4_22),
.matrixC4_23(matrixC4_23),
.matrixC4_24(matrixC4_24),
.matrixC4_25(matrixC4_25),
.matrixC4_26(matrixC4_26),
.matrixC4_27(matrixC4_27),
.matrixC4_28(matrixC4_28),
.matrixC4_29(matrixC4_29),
.matrixC4_30(matrixC4_30),
.matrixC4_31(matrixC4_31),
.matrixC5_0(matrixC5_0),
.matrixC5_1(matrixC5_1),
.matrixC5_2(matrixC5_2),
.matrixC5_3(matrixC5_3),
.matrixC5_4(matrixC5_4),
.matrixC5_5(matrixC5_5),
.matrixC5_6(matrixC5_6),
.matrixC5_7(matrixC5_7),
.matrixC5_8(matrixC5_8),
.matrixC5_9(matrixC5_9),
.matrixC5_10(matrixC5_10),
.matrixC5_11(matrixC5_11),
.matrixC5_12(matrixC5_12),
.matrixC5_13(matrixC5_13),
.matrixC5_14(matrixC5_14),
.matrixC5_15(matrixC5_15),
.matrixC5_16(matrixC5_16),
.matrixC5_17(matrixC5_17),
.matrixC5_18(matrixC5_18),
.matrixC5_19(matrixC5_19),
.matrixC5_20(matrixC5_20),
.matrixC5_21(matrixC5_21),
.matrixC5_22(matrixC5_22),
.matrixC5_23(matrixC5_23),
.matrixC5_24(matrixC5_24),
.matrixC5_25(matrixC5_25),
.matrixC5_26(matrixC5_26),
.matrixC5_27(matrixC5_27),
.matrixC5_28(matrixC5_28),
.matrixC5_29(matrixC5_29),
.matrixC5_30(matrixC5_30),
.matrixC5_31(matrixC5_31),
.matrixC6_0(matrixC6_0),
.matrixC6_1(matrixC6_1),
.matrixC6_2(matrixC6_2),
.matrixC6_3(matrixC6_3),
.matrixC6_4(matrixC6_4),
.matrixC6_5(matrixC6_5),
.matrixC6_6(matrixC6_6),
.matrixC6_7(matrixC6_7),
.matrixC6_8(matrixC6_8),
.matrixC6_9(matrixC6_9),
.matrixC6_10(matrixC6_10),
.matrixC6_11(matrixC6_11),
.matrixC6_12(matrixC6_12),
.matrixC6_13(matrixC6_13),
.matrixC6_14(matrixC6_14),
.matrixC6_15(matrixC6_15),
.matrixC6_16(matrixC6_16),
.matrixC6_17(matrixC6_17),
.matrixC6_18(matrixC6_18),
.matrixC6_19(matrixC6_19),
.matrixC6_20(matrixC6_20),
.matrixC6_21(matrixC6_21),
.matrixC6_22(matrixC6_22),
.matrixC6_23(matrixC6_23),
.matrixC6_24(matrixC6_24),
.matrixC6_25(matrixC6_25),
.matrixC6_26(matrixC6_26),
.matrixC6_27(matrixC6_27),
.matrixC6_28(matrixC6_28),
.matrixC6_29(matrixC6_29),
.matrixC6_30(matrixC6_30),
.matrixC6_31(matrixC6_31),
.matrixC7_0(matrixC7_0),
.matrixC7_1(matrixC7_1),
.matrixC7_2(matrixC7_2),
.matrixC7_3(matrixC7_3),
.matrixC7_4(matrixC7_4),
.matrixC7_5(matrixC7_5),
.matrixC7_6(matrixC7_6),
.matrixC7_7(matrixC7_7),
.matrixC7_8(matrixC7_8),
.matrixC7_9(matrixC7_9),
.matrixC7_10(matrixC7_10),
.matrixC7_11(matrixC7_11),
.matrixC7_12(matrixC7_12),
.matrixC7_13(matrixC7_13),
.matrixC7_14(matrixC7_14),
.matrixC7_15(matrixC7_15),
.matrixC7_16(matrixC7_16),
.matrixC7_17(matrixC7_17),
.matrixC7_18(matrixC7_18),
.matrixC7_19(matrixC7_19),
.matrixC7_20(matrixC7_20),
.matrixC7_21(matrixC7_21),
.matrixC7_22(matrixC7_22),
.matrixC7_23(matrixC7_23),
.matrixC7_24(matrixC7_24),
.matrixC7_25(matrixC7_25),
.matrixC7_26(matrixC7_26),
.matrixC7_27(matrixC7_27),
.matrixC7_28(matrixC7_28),
.matrixC7_29(matrixC7_29),
.matrixC7_30(matrixC7_30),
.matrixC7_31(matrixC7_31),
.matrixC8_0(matrixC8_0),
.matrixC8_1(matrixC8_1),
.matrixC8_2(matrixC8_2),
.matrixC8_3(matrixC8_3),
.matrixC8_4(matrixC8_4),
.matrixC8_5(matrixC8_5),
.matrixC8_6(matrixC8_6),
.matrixC8_7(matrixC8_7),
.matrixC8_8(matrixC8_8),
.matrixC8_9(matrixC8_9),
.matrixC8_10(matrixC8_10),
.matrixC8_11(matrixC8_11),
.matrixC8_12(matrixC8_12),
.matrixC8_13(matrixC8_13),
.matrixC8_14(matrixC8_14),
.matrixC8_15(matrixC8_15),
.matrixC8_16(matrixC8_16),
.matrixC8_17(matrixC8_17),
.matrixC8_18(matrixC8_18),
.matrixC8_19(matrixC8_19),
.matrixC8_20(matrixC8_20),
.matrixC8_21(matrixC8_21),
.matrixC8_22(matrixC8_22),
.matrixC8_23(matrixC8_23),
.matrixC8_24(matrixC8_24),
.matrixC8_25(matrixC8_25),
.matrixC8_26(matrixC8_26),
.matrixC8_27(matrixC8_27),
.matrixC8_28(matrixC8_28),
.matrixC8_29(matrixC8_29),
.matrixC8_30(matrixC8_30),
.matrixC8_31(matrixC8_31),
.matrixC9_0(matrixC9_0),
.matrixC9_1(matrixC9_1),
.matrixC9_2(matrixC9_2),
.matrixC9_3(matrixC9_3),
.matrixC9_4(matrixC9_4),
.matrixC9_5(matrixC9_5),
.matrixC9_6(matrixC9_6),
.matrixC9_7(matrixC9_7),
.matrixC9_8(matrixC9_8),
.matrixC9_9(matrixC9_9),
.matrixC9_10(matrixC9_10),
.matrixC9_11(matrixC9_11),
.matrixC9_12(matrixC9_12),
.matrixC9_13(matrixC9_13),
.matrixC9_14(matrixC9_14),
.matrixC9_15(matrixC9_15),
.matrixC9_16(matrixC9_16),
.matrixC9_17(matrixC9_17),
.matrixC9_18(matrixC9_18),
.matrixC9_19(matrixC9_19),
.matrixC9_20(matrixC9_20),
.matrixC9_21(matrixC9_21),
.matrixC9_22(matrixC9_22),
.matrixC9_23(matrixC9_23),
.matrixC9_24(matrixC9_24),
.matrixC9_25(matrixC9_25),
.matrixC9_26(matrixC9_26),
.matrixC9_27(matrixC9_27),
.matrixC9_28(matrixC9_28),
.matrixC9_29(matrixC9_29),
.matrixC9_30(matrixC9_30),
.matrixC9_31(matrixC9_31),
.matrixC10_0(matrixC10_0),
.matrixC10_1(matrixC10_1),
.matrixC10_2(matrixC10_2),
.matrixC10_3(matrixC10_3),
.matrixC10_4(matrixC10_4),
.matrixC10_5(matrixC10_5),
.matrixC10_6(matrixC10_6),
.matrixC10_7(matrixC10_7),
.matrixC10_8(matrixC10_8),
.matrixC10_9(matrixC10_9),
.matrixC10_10(matrixC10_10),
.matrixC10_11(matrixC10_11),
.matrixC10_12(matrixC10_12),
.matrixC10_13(matrixC10_13),
.matrixC10_14(matrixC10_14),
.matrixC10_15(matrixC10_15),
.matrixC10_16(matrixC10_16),
.matrixC10_17(matrixC10_17),
.matrixC10_18(matrixC10_18),
.matrixC10_19(matrixC10_19),
.matrixC10_20(matrixC10_20),
.matrixC10_21(matrixC10_21),
.matrixC10_22(matrixC10_22),
.matrixC10_23(matrixC10_23),
.matrixC10_24(matrixC10_24),
.matrixC10_25(matrixC10_25),
.matrixC10_26(matrixC10_26),
.matrixC10_27(matrixC10_27),
.matrixC10_28(matrixC10_28),
.matrixC10_29(matrixC10_29),
.matrixC10_30(matrixC10_30),
.matrixC10_31(matrixC10_31),
.matrixC11_0(matrixC11_0),
.matrixC11_1(matrixC11_1),
.matrixC11_2(matrixC11_2),
.matrixC11_3(matrixC11_3),
.matrixC11_4(matrixC11_4),
.matrixC11_5(matrixC11_5),
.matrixC11_6(matrixC11_6),
.matrixC11_7(matrixC11_7),
.matrixC11_8(matrixC11_8),
.matrixC11_9(matrixC11_9),
.matrixC11_10(matrixC11_10),
.matrixC11_11(matrixC11_11),
.matrixC11_12(matrixC11_12),
.matrixC11_13(matrixC11_13),
.matrixC11_14(matrixC11_14),
.matrixC11_15(matrixC11_15),
.matrixC11_16(matrixC11_16),
.matrixC11_17(matrixC11_17),
.matrixC11_18(matrixC11_18),
.matrixC11_19(matrixC11_19),
.matrixC11_20(matrixC11_20),
.matrixC11_21(matrixC11_21),
.matrixC11_22(matrixC11_22),
.matrixC11_23(matrixC11_23),
.matrixC11_24(matrixC11_24),
.matrixC11_25(matrixC11_25),
.matrixC11_26(matrixC11_26),
.matrixC11_27(matrixC11_27),
.matrixC11_28(matrixC11_28),
.matrixC11_29(matrixC11_29),
.matrixC11_30(matrixC11_30),
.matrixC11_31(matrixC11_31),
.matrixC12_0(matrixC12_0),
.matrixC12_1(matrixC12_1),
.matrixC12_2(matrixC12_2),
.matrixC12_3(matrixC12_3),
.matrixC12_4(matrixC12_4),
.matrixC12_5(matrixC12_5),
.matrixC12_6(matrixC12_6),
.matrixC12_7(matrixC12_7),
.matrixC12_8(matrixC12_8),
.matrixC12_9(matrixC12_9),
.matrixC12_10(matrixC12_10),
.matrixC12_11(matrixC12_11),
.matrixC12_12(matrixC12_12),
.matrixC12_13(matrixC12_13),
.matrixC12_14(matrixC12_14),
.matrixC12_15(matrixC12_15),
.matrixC12_16(matrixC12_16),
.matrixC12_17(matrixC12_17),
.matrixC12_18(matrixC12_18),
.matrixC12_19(matrixC12_19),
.matrixC12_20(matrixC12_20),
.matrixC12_21(matrixC12_21),
.matrixC12_22(matrixC12_22),
.matrixC12_23(matrixC12_23),
.matrixC12_24(matrixC12_24),
.matrixC12_25(matrixC12_25),
.matrixC12_26(matrixC12_26),
.matrixC12_27(matrixC12_27),
.matrixC12_28(matrixC12_28),
.matrixC12_29(matrixC12_29),
.matrixC12_30(matrixC12_30),
.matrixC12_31(matrixC12_31),
.matrixC13_0(matrixC13_0),
.matrixC13_1(matrixC13_1),
.matrixC13_2(matrixC13_2),
.matrixC13_3(matrixC13_3),
.matrixC13_4(matrixC13_4),
.matrixC13_5(matrixC13_5),
.matrixC13_6(matrixC13_6),
.matrixC13_7(matrixC13_7),
.matrixC13_8(matrixC13_8),
.matrixC13_9(matrixC13_9),
.matrixC13_10(matrixC13_10),
.matrixC13_11(matrixC13_11),
.matrixC13_12(matrixC13_12),
.matrixC13_13(matrixC13_13),
.matrixC13_14(matrixC13_14),
.matrixC13_15(matrixC13_15),
.matrixC13_16(matrixC13_16),
.matrixC13_17(matrixC13_17),
.matrixC13_18(matrixC13_18),
.matrixC13_19(matrixC13_19),
.matrixC13_20(matrixC13_20),
.matrixC13_21(matrixC13_21),
.matrixC13_22(matrixC13_22),
.matrixC13_23(matrixC13_23),
.matrixC13_24(matrixC13_24),
.matrixC13_25(matrixC13_25),
.matrixC13_26(matrixC13_26),
.matrixC13_27(matrixC13_27),
.matrixC13_28(matrixC13_28),
.matrixC13_29(matrixC13_29),
.matrixC13_30(matrixC13_30),
.matrixC13_31(matrixC13_31),
.matrixC14_0(matrixC14_0),
.matrixC14_1(matrixC14_1),
.matrixC14_2(matrixC14_2),
.matrixC14_3(matrixC14_3),
.matrixC14_4(matrixC14_4),
.matrixC14_5(matrixC14_5),
.matrixC14_6(matrixC14_6),
.matrixC14_7(matrixC14_7),
.matrixC14_8(matrixC14_8),
.matrixC14_9(matrixC14_9),
.matrixC14_10(matrixC14_10),
.matrixC14_11(matrixC14_11),
.matrixC14_12(matrixC14_12),
.matrixC14_13(matrixC14_13),
.matrixC14_14(matrixC14_14),
.matrixC14_15(matrixC14_15),
.matrixC14_16(matrixC14_16),
.matrixC14_17(matrixC14_17),
.matrixC14_18(matrixC14_18),
.matrixC14_19(matrixC14_19),
.matrixC14_20(matrixC14_20),
.matrixC14_21(matrixC14_21),
.matrixC14_22(matrixC14_22),
.matrixC14_23(matrixC14_23),
.matrixC14_24(matrixC14_24),
.matrixC14_25(matrixC14_25),
.matrixC14_26(matrixC14_26),
.matrixC14_27(matrixC14_27),
.matrixC14_28(matrixC14_28),
.matrixC14_29(matrixC14_29),
.matrixC14_30(matrixC14_30),
.matrixC14_31(matrixC14_31),
.matrixC15_0(matrixC15_0),
.matrixC15_1(matrixC15_1),
.matrixC15_2(matrixC15_2),
.matrixC15_3(matrixC15_3),
.matrixC15_4(matrixC15_4),
.matrixC15_5(matrixC15_5),
.matrixC15_6(matrixC15_6),
.matrixC15_7(matrixC15_7),
.matrixC15_8(matrixC15_8),
.matrixC15_9(matrixC15_9),
.matrixC15_10(matrixC15_10),
.matrixC15_11(matrixC15_11),
.matrixC15_12(matrixC15_12),
.matrixC15_13(matrixC15_13),
.matrixC15_14(matrixC15_14),
.matrixC15_15(matrixC15_15),
.matrixC15_16(matrixC15_16),
.matrixC15_17(matrixC15_17),
.matrixC15_18(matrixC15_18),
.matrixC15_19(matrixC15_19),
.matrixC15_20(matrixC15_20),
.matrixC15_21(matrixC15_21),
.matrixC15_22(matrixC15_22),
.matrixC15_23(matrixC15_23),
.matrixC15_24(matrixC15_24),
.matrixC15_25(matrixC15_25),
.matrixC15_26(matrixC15_26),
.matrixC15_27(matrixC15_27),
.matrixC15_28(matrixC15_28),
.matrixC15_29(matrixC15_29),
.matrixC15_30(matrixC15_30),
.matrixC15_31(matrixC15_31),
.matrixC16_0(matrixC16_0),
.matrixC16_1(matrixC16_1),
.matrixC16_2(matrixC16_2),
.matrixC16_3(matrixC16_3),
.matrixC16_4(matrixC16_4),
.matrixC16_5(matrixC16_5),
.matrixC16_6(matrixC16_6),
.matrixC16_7(matrixC16_7),
.matrixC16_8(matrixC16_8),
.matrixC16_9(matrixC16_9),
.matrixC16_10(matrixC16_10),
.matrixC16_11(matrixC16_11),
.matrixC16_12(matrixC16_12),
.matrixC16_13(matrixC16_13),
.matrixC16_14(matrixC16_14),
.matrixC16_15(matrixC16_15),
.matrixC16_16(matrixC16_16),
.matrixC16_17(matrixC16_17),
.matrixC16_18(matrixC16_18),
.matrixC16_19(matrixC16_19),
.matrixC16_20(matrixC16_20),
.matrixC16_21(matrixC16_21),
.matrixC16_22(matrixC16_22),
.matrixC16_23(matrixC16_23),
.matrixC16_24(matrixC16_24),
.matrixC16_25(matrixC16_25),
.matrixC16_26(matrixC16_26),
.matrixC16_27(matrixC16_27),
.matrixC16_28(matrixC16_28),
.matrixC16_29(matrixC16_29),
.matrixC16_30(matrixC16_30),
.matrixC16_31(matrixC16_31),
.matrixC17_0(matrixC17_0),
.matrixC17_1(matrixC17_1),
.matrixC17_2(matrixC17_2),
.matrixC17_3(matrixC17_3),
.matrixC17_4(matrixC17_4),
.matrixC17_5(matrixC17_5),
.matrixC17_6(matrixC17_6),
.matrixC17_7(matrixC17_7),
.matrixC17_8(matrixC17_8),
.matrixC17_9(matrixC17_9),
.matrixC17_10(matrixC17_10),
.matrixC17_11(matrixC17_11),
.matrixC17_12(matrixC17_12),
.matrixC17_13(matrixC17_13),
.matrixC17_14(matrixC17_14),
.matrixC17_15(matrixC17_15),
.matrixC17_16(matrixC17_16),
.matrixC17_17(matrixC17_17),
.matrixC17_18(matrixC17_18),
.matrixC17_19(matrixC17_19),
.matrixC17_20(matrixC17_20),
.matrixC17_21(matrixC17_21),
.matrixC17_22(matrixC17_22),
.matrixC17_23(matrixC17_23),
.matrixC17_24(matrixC17_24),
.matrixC17_25(matrixC17_25),
.matrixC17_26(matrixC17_26),
.matrixC17_27(matrixC17_27),
.matrixC17_28(matrixC17_28),
.matrixC17_29(matrixC17_29),
.matrixC17_30(matrixC17_30),
.matrixC17_31(matrixC17_31),
.matrixC18_0(matrixC18_0),
.matrixC18_1(matrixC18_1),
.matrixC18_2(matrixC18_2),
.matrixC18_3(matrixC18_3),
.matrixC18_4(matrixC18_4),
.matrixC18_5(matrixC18_5),
.matrixC18_6(matrixC18_6),
.matrixC18_7(matrixC18_7),
.matrixC18_8(matrixC18_8),
.matrixC18_9(matrixC18_9),
.matrixC18_10(matrixC18_10),
.matrixC18_11(matrixC18_11),
.matrixC18_12(matrixC18_12),
.matrixC18_13(matrixC18_13),
.matrixC18_14(matrixC18_14),
.matrixC18_15(matrixC18_15),
.matrixC18_16(matrixC18_16),
.matrixC18_17(matrixC18_17),
.matrixC18_18(matrixC18_18),
.matrixC18_19(matrixC18_19),
.matrixC18_20(matrixC18_20),
.matrixC18_21(matrixC18_21),
.matrixC18_22(matrixC18_22),
.matrixC18_23(matrixC18_23),
.matrixC18_24(matrixC18_24),
.matrixC18_25(matrixC18_25),
.matrixC18_26(matrixC18_26),
.matrixC18_27(matrixC18_27),
.matrixC18_28(matrixC18_28),
.matrixC18_29(matrixC18_29),
.matrixC18_30(matrixC18_30),
.matrixC18_31(matrixC18_31),
.matrixC19_0(matrixC19_0),
.matrixC19_1(matrixC19_1),
.matrixC19_2(matrixC19_2),
.matrixC19_3(matrixC19_3),
.matrixC19_4(matrixC19_4),
.matrixC19_5(matrixC19_5),
.matrixC19_6(matrixC19_6),
.matrixC19_7(matrixC19_7),
.matrixC19_8(matrixC19_8),
.matrixC19_9(matrixC19_9),
.matrixC19_10(matrixC19_10),
.matrixC19_11(matrixC19_11),
.matrixC19_12(matrixC19_12),
.matrixC19_13(matrixC19_13),
.matrixC19_14(matrixC19_14),
.matrixC19_15(matrixC19_15),
.matrixC19_16(matrixC19_16),
.matrixC19_17(matrixC19_17),
.matrixC19_18(matrixC19_18),
.matrixC19_19(matrixC19_19),
.matrixC19_20(matrixC19_20),
.matrixC19_21(matrixC19_21),
.matrixC19_22(matrixC19_22),
.matrixC19_23(matrixC19_23),
.matrixC19_24(matrixC19_24),
.matrixC19_25(matrixC19_25),
.matrixC19_26(matrixC19_26),
.matrixC19_27(matrixC19_27),
.matrixC19_28(matrixC19_28),
.matrixC19_29(matrixC19_29),
.matrixC19_30(matrixC19_30),
.matrixC19_31(matrixC19_31),
.matrixC20_0(matrixC20_0),
.matrixC20_1(matrixC20_1),
.matrixC20_2(matrixC20_2),
.matrixC20_3(matrixC20_3),
.matrixC20_4(matrixC20_4),
.matrixC20_5(matrixC20_5),
.matrixC20_6(matrixC20_6),
.matrixC20_7(matrixC20_7),
.matrixC20_8(matrixC20_8),
.matrixC20_9(matrixC20_9),
.matrixC20_10(matrixC20_10),
.matrixC20_11(matrixC20_11),
.matrixC20_12(matrixC20_12),
.matrixC20_13(matrixC20_13),
.matrixC20_14(matrixC20_14),
.matrixC20_15(matrixC20_15),
.matrixC20_16(matrixC20_16),
.matrixC20_17(matrixC20_17),
.matrixC20_18(matrixC20_18),
.matrixC20_19(matrixC20_19),
.matrixC20_20(matrixC20_20),
.matrixC20_21(matrixC20_21),
.matrixC20_22(matrixC20_22),
.matrixC20_23(matrixC20_23),
.matrixC20_24(matrixC20_24),
.matrixC20_25(matrixC20_25),
.matrixC20_26(matrixC20_26),
.matrixC20_27(matrixC20_27),
.matrixC20_28(matrixC20_28),
.matrixC20_29(matrixC20_29),
.matrixC20_30(matrixC20_30),
.matrixC20_31(matrixC20_31),
.matrixC21_0(matrixC21_0),
.matrixC21_1(matrixC21_1),
.matrixC21_2(matrixC21_2),
.matrixC21_3(matrixC21_3),
.matrixC21_4(matrixC21_4),
.matrixC21_5(matrixC21_5),
.matrixC21_6(matrixC21_6),
.matrixC21_7(matrixC21_7),
.matrixC21_8(matrixC21_8),
.matrixC21_9(matrixC21_9),
.matrixC21_10(matrixC21_10),
.matrixC21_11(matrixC21_11),
.matrixC21_12(matrixC21_12),
.matrixC21_13(matrixC21_13),
.matrixC21_14(matrixC21_14),
.matrixC21_15(matrixC21_15),
.matrixC21_16(matrixC21_16),
.matrixC21_17(matrixC21_17),
.matrixC21_18(matrixC21_18),
.matrixC21_19(matrixC21_19),
.matrixC21_20(matrixC21_20),
.matrixC21_21(matrixC21_21),
.matrixC21_22(matrixC21_22),
.matrixC21_23(matrixC21_23),
.matrixC21_24(matrixC21_24),
.matrixC21_25(matrixC21_25),
.matrixC21_26(matrixC21_26),
.matrixC21_27(matrixC21_27),
.matrixC21_28(matrixC21_28),
.matrixC21_29(matrixC21_29),
.matrixC21_30(matrixC21_30),
.matrixC21_31(matrixC21_31),
.matrixC22_0(matrixC22_0),
.matrixC22_1(matrixC22_1),
.matrixC22_2(matrixC22_2),
.matrixC22_3(matrixC22_3),
.matrixC22_4(matrixC22_4),
.matrixC22_5(matrixC22_5),
.matrixC22_6(matrixC22_6),
.matrixC22_7(matrixC22_7),
.matrixC22_8(matrixC22_8),
.matrixC22_9(matrixC22_9),
.matrixC22_10(matrixC22_10),
.matrixC22_11(matrixC22_11),
.matrixC22_12(matrixC22_12),
.matrixC22_13(matrixC22_13),
.matrixC22_14(matrixC22_14),
.matrixC22_15(matrixC22_15),
.matrixC22_16(matrixC22_16),
.matrixC22_17(matrixC22_17),
.matrixC22_18(matrixC22_18),
.matrixC22_19(matrixC22_19),
.matrixC22_20(matrixC22_20),
.matrixC22_21(matrixC22_21),
.matrixC22_22(matrixC22_22),
.matrixC22_23(matrixC22_23),
.matrixC22_24(matrixC22_24),
.matrixC22_25(matrixC22_25),
.matrixC22_26(matrixC22_26),
.matrixC22_27(matrixC22_27),
.matrixC22_28(matrixC22_28),
.matrixC22_29(matrixC22_29),
.matrixC22_30(matrixC22_30),
.matrixC22_31(matrixC22_31),
.matrixC23_0(matrixC23_0),
.matrixC23_1(matrixC23_1),
.matrixC23_2(matrixC23_2),
.matrixC23_3(matrixC23_3),
.matrixC23_4(matrixC23_4),
.matrixC23_5(matrixC23_5),
.matrixC23_6(matrixC23_6),
.matrixC23_7(matrixC23_7),
.matrixC23_8(matrixC23_8),
.matrixC23_9(matrixC23_9),
.matrixC23_10(matrixC23_10),
.matrixC23_11(matrixC23_11),
.matrixC23_12(matrixC23_12),
.matrixC23_13(matrixC23_13),
.matrixC23_14(matrixC23_14),
.matrixC23_15(matrixC23_15),
.matrixC23_16(matrixC23_16),
.matrixC23_17(matrixC23_17),
.matrixC23_18(matrixC23_18),
.matrixC23_19(matrixC23_19),
.matrixC23_20(matrixC23_20),
.matrixC23_21(matrixC23_21),
.matrixC23_22(matrixC23_22),
.matrixC23_23(matrixC23_23),
.matrixC23_24(matrixC23_24),
.matrixC23_25(matrixC23_25),
.matrixC23_26(matrixC23_26),
.matrixC23_27(matrixC23_27),
.matrixC23_28(matrixC23_28),
.matrixC23_29(matrixC23_29),
.matrixC23_30(matrixC23_30),
.matrixC23_31(matrixC23_31),
.matrixC24_0(matrixC24_0),
.matrixC24_1(matrixC24_1),
.matrixC24_2(matrixC24_2),
.matrixC24_3(matrixC24_3),
.matrixC24_4(matrixC24_4),
.matrixC24_5(matrixC24_5),
.matrixC24_6(matrixC24_6),
.matrixC24_7(matrixC24_7),
.matrixC24_8(matrixC24_8),
.matrixC24_9(matrixC24_9),
.matrixC24_10(matrixC24_10),
.matrixC24_11(matrixC24_11),
.matrixC24_12(matrixC24_12),
.matrixC24_13(matrixC24_13),
.matrixC24_14(matrixC24_14),
.matrixC24_15(matrixC24_15),
.matrixC24_16(matrixC24_16),
.matrixC24_17(matrixC24_17),
.matrixC24_18(matrixC24_18),
.matrixC24_19(matrixC24_19),
.matrixC24_20(matrixC24_20),
.matrixC24_21(matrixC24_21),
.matrixC24_22(matrixC24_22),
.matrixC24_23(matrixC24_23),
.matrixC24_24(matrixC24_24),
.matrixC24_25(matrixC24_25),
.matrixC24_26(matrixC24_26),
.matrixC24_27(matrixC24_27),
.matrixC24_28(matrixC24_28),
.matrixC24_29(matrixC24_29),
.matrixC24_30(matrixC24_30),
.matrixC24_31(matrixC24_31),
.matrixC25_0(matrixC25_0),
.matrixC25_1(matrixC25_1),
.matrixC25_2(matrixC25_2),
.matrixC25_3(matrixC25_3),
.matrixC25_4(matrixC25_4),
.matrixC25_5(matrixC25_5),
.matrixC25_6(matrixC25_6),
.matrixC25_7(matrixC25_7),
.matrixC25_8(matrixC25_8),
.matrixC25_9(matrixC25_9),
.matrixC25_10(matrixC25_10),
.matrixC25_11(matrixC25_11),
.matrixC25_12(matrixC25_12),
.matrixC25_13(matrixC25_13),
.matrixC25_14(matrixC25_14),
.matrixC25_15(matrixC25_15),
.matrixC25_16(matrixC25_16),
.matrixC25_17(matrixC25_17),
.matrixC25_18(matrixC25_18),
.matrixC25_19(matrixC25_19),
.matrixC25_20(matrixC25_20),
.matrixC25_21(matrixC25_21),
.matrixC25_22(matrixC25_22),
.matrixC25_23(matrixC25_23),
.matrixC25_24(matrixC25_24),
.matrixC25_25(matrixC25_25),
.matrixC25_26(matrixC25_26),
.matrixC25_27(matrixC25_27),
.matrixC25_28(matrixC25_28),
.matrixC25_29(matrixC25_29),
.matrixC25_30(matrixC25_30),
.matrixC25_31(matrixC25_31),
.matrixC26_0(matrixC26_0),
.matrixC26_1(matrixC26_1),
.matrixC26_2(matrixC26_2),
.matrixC26_3(matrixC26_3),
.matrixC26_4(matrixC26_4),
.matrixC26_5(matrixC26_5),
.matrixC26_6(matrixC26_6),
.matrixC26_7(matrixC26_7),
.matrixC26_8(matrixC26_8),
.matrixC26_9(matrixC26_9),
.matrixC26_10(matrixC26_10),
.matrixC26_11(matrixC26_11),
.matrixC26_12(matrixC26_12),
.matrixC26_13(matrixC26_13),
.matrixC26_14(matrixC26_14),
.matrixC26_15(matrixC26_15),
.matrixC26_16(matrixC26_16),
.matrixC26_17(matrixC26_17),
.matrixC26_18(matrixC26_18),
.matrixC26_19(matrixC26_19),
.matrixC26_20(matrixC26_20),
.matrixC26_21(matrixC26_21),
.matrixC26_22(matrixC26_22),
.matrixC26_23(matrixC26_23),
.matrixC26_24(matrixC26_24),
.matrixC26_25(matrixC26_25),
.matrixC26_26(matrixC26_26),
.matrixC26_27(matrixC26_27),
.matrixC26_28(matrixC26_28),
.matrixC26_29(matrixC26_29),
.matrixC26_30(matrixC26_30),
.matrixC26_31(matrixC26_31),
.matrixC27_0(matrixC27_0),
.matrixC27_1(matrixC27_1),
.matrixC27_2(matrixC27_2),
.matrixC27_3(matrixC27_3),
.matrixC27_4(matrixC27_4),
.matrixC27_5(matrixC27_5),
.matrixC27_6(matrixC27_6),
.matrixC27_7(matrixC27_7),
.matrixC27_8(matrixC27_8),
.matrixC27_9(matrixC27_9),
.matrixC27_10(matrixC27_10),
.matrixC27_11(matrixC27_11),
.matrixC27_12(matrixC27_12),
.matrixC27_13(matrixC27_13),
.matrixC27_14(matrixC27_14),
.matrixC27_15(matrixC27_15),
.matrixC27_16(matrixC27_16),
.matrixC27_17(matrixC27_17),
.matrixC27_18(matrixC27_18),
.matrixC27_19(matrixC27_19),
.matrixC27_20(matrixC27_20),
.matrixC27_21(matrixC27_21),
.matrixC27_22(matrixC27_22),
.matrixC27_23(matrixC27_23),
.matrixC27_24(matrixC27_24),
.matrixC27_25(matrixC27_25),
.matrixC27_26(matrixC27_26),
.matrixC27_27(matrixC27_27),
.matrixC27_28(matrixC27_28),
.matrixC27_29(matrixC27_29),
.matrixC27_30(matrixC27_30),
.matrixC27_31(matrixC27_31),
.matrixC28_0(matrixC28_0),
.matrixC28_1(matrixC28_1),
.matrixC28_2(matrixC28_2),
.matrixC28_3(matrixC28_3),
.matrixC28_4(matrixC28_4),
.matrixC28_5(matrixC28_5),
.matrixC28_6(matrixC28_6),
.matrixC28_7(matrixC28_7),
.matrixC28_8(matrixC28_8),
.matrixC28_9(matrixC28_9),
.matrixC28_10(matrixC28_10),
.matrixC28_11(matrixC28_11),
.matrixC28_12(matrixC28_12),
.matrixC28_13(matrixC28_13),
.matrixC28_14(matrixC28_14),
.matrixC28_15(matrixC28_15),
.matrixC28_16(matrixC28_16),
.matrixC28_17(matrixC28_17),
.matrixC28_18(matrixC28_18),
.matrixC28_19(matrixC28_19),
.matrixC28_20(matrixC28_20),
.matrixC28_21(matrixC28_21),
.matrixC28_22(matrixC28_22),
.matrixC28_23(matrixC28_23),
.matrixC28_24(matrixC28_24),
.matrixC28_25(matrixC28_25),
.matrixC28_26(matrixC28_26),
.matrixC28_27(matrixC28_27),
.matrixC28_28(matrixC28_28),
.matrixC28_29(matrixC28_29),
.matrixC28_30(matrixC28_30),
.matrixC28_31(matrixC28_31),
.matrixC29_0(matrixC29_0),
.matrixC29_1(matrixC29_1),
.matrixC29_2(matrixC29_2),
.matrixC29_3(matrixC29_3),
.matrixC29_4(matrixC29_4),
.matrixC29_5(matrixC29_5),
.matrixC29_6(matrixC29_6),
.matrixC29_7(matrixC29_7),
.matrixC29_8(matrixC29_8),
.matrixC29_9(matrixC29_9),
.matrixC29_10(matrixC29_10),
.matrixC29_11(matrixC29_11),
.matrixC29_12(matrixC29_12),
.matrixC29_13(matrixC29_13),
.matrixC29_14(matrixC29_14),
.matrixC29_15(matrixC29_15),
.matrixC29_16(matrixC29_16),
.matrixC29_17(matrixC29_17),
.matrixC29_18(matrixC29_18),
.matrixC29_19(matrixC29_19),
.matrixC29_20(matrixC29_20),
.matrixC29_21(matrixC29_21),
.matrixC29_22(matrixC29_22),
.matrixC29_23(matrixC29_23),
.matrixC29_24(matrixC29_24),
.matrixC29_25(matrixC29_25),
.matrixC29_26(matrixC29_26),
.matrixC29_27(matrixC29_27),
.matrixC29_28(matrixC29_28),
.matrixC29_29(matrixC29_29),
.matrixC29_30(matrixC29_30),
.matrixC29_31(matrixC29_31),
.matrixC30_0(matrixC30_0),
.matrixC30_1(matrixC30_1),
.matrixC30_2(matrixC30_2),
.matrixC30_3(matrixC30_3),
.matrixC30_4(matrixC30_4),
.matrixC30_5(matrixC30_5),
.matrixC30_6(matrixC30_6),
.matrixC30_7(matrixC30_7),
.matrixC30_8(matrixC30_8),
.matrixC30_9(matrixC30_9),
.matrixC30_10(matrixC30_10),
.matrixC30_11(matrixC30_11),
.matrixC30_12(matrixC30_12),
.matrixC30_13(matrixC30_13),
.matrixC30_14(matrixC30_14),
.matrixC30_15(matrixC30_15),
.matrixC30_16(matrixC30_16),
.matrixC30_17(matrixC30_17),
.matrixC30_18(matrixC30_18),
.matrixC30_19(matrixC30_19),
.matrixC30_20(matrixC30_20),
.matrixC30_21(matrixC30_21),
.matrixC30_22(matrixC30_22),
.matrixC30_23(matrixC30_23),
.matrixC30_24(matrixC30_24),
.matrixC30_25(matrixC30_25),
.matrixC30_26(matrixC30_26),
.matrixC30_27(matrixC30_27),
.matrixC30_28(matrixC30_28),
.matrixC30_29(matrixC30_29),
.matrixC30_30(matrixC30_30),
.matrixC30_31(matrixC30_31),
.matrixC31_0(matrixC31_0),
.matrixC31_1(matrixC31_1),
.matrixC31_2(matrixC31_2),
.matrixC31_3(matrixC31_3),
.matrixC31_4(matrixC31_4),
.matrixC31_5(matrixC31_5),
.matrixC31_6(matrixC31_6),
.matrixC31_7(matrixC31_7),
.matrixC31_8(matrixC31_8),
.matrixC31_9(matrixC31_9),
.matrixC31_10(matrixC31_10),
.matrixC31_11(matrixC31_11),
.matrixC31_12(matrixC31_12),
.matrixC31_13(matrixC31_13),
.matrixC31_14(matrixC31_14),
.matrixC31_15(matrixC31_15),
.matrixC31_16(matrixC31_16),
.matrixC31_17(matrixC31_17),
.matrixC31_18(matrixC31_18),
.matrixC31_19(matrixC31_19),
.matrixC31_20(matrixC31_20),
.matrixC31_21(matrixC31_21),
.matrixC31_22(matrixC31_22),
.matrixC31_23(matrixC31_23),
.matrixC31_24(matrixC31_24),
.matrixC31_25(matrixC31_25),
.matrixC31_26(matrixC31_26),
.matrixC31_27(matrixC31_27),
.matrixC31_28(matrixC31_28),
.matrixC31_29(matrixC31_29),
.matrixC31_30(matrixC31_30),
.matrixC31_31(matrixC31_31),

.clk(clk),
.reset(reset)
);

//////////////////////////////////////////////////////////////////////////
// Instantiations of the actual PEs
//////////////////////////////////////////////////////////////////////////
systolic_pe_matrix u_systolic_pe_matrix(
.clk(clk),
.reset(reset),
.pe_reset(pe_reset),
.start_mat_mul(start_mat_mul),
.a0(a0),
.a1(a1),
.a2(a2),
.a3(a3),
.a4(a4),
.a5(a5),
.a6(a6),
.a7(a7),
.a8(a8),
.a9(a9),
.a10(a10),
.a11(a11),
.a12(a12),
.a13(a13),
.a14(a14),
.a15(a15),
.a16(a16),
.a17(a17),
.a18(a18),
.a19(a19),
.a20(a20),
.a21(a21),
.a22(a22),
.a23(a23),
.a24(a24),
.a25(a25),
.a26(a26),
.a27(a27),
.a28(a28),
.a29(a29),
.a30(a30),
.a31(a31),
.b0(b0),
.b1(b1),
.b2(b2),
.b3(b3),
.b4(b4),
.b5(b5),
.b6(b6),
.b7(b7),
.b8(b8),
.b9(b9),
.b10(b10),
.b11(b11),
.b12(b12),
.b13(b13),
.b14(b14),
.b15(b15),
.b16(b16),
.b17(b17),
.b18(b18),
.b19(b19),
.b20(b20),
.b21(b21),
.b22(b22),
.b23(b23),
.b24(b24),
.b25(b25),
.b26(b26),
.b27(b27),
.b28(b28),
.b29(b29),
.b30(b30),
.b31(b31),
.matrixC0_0(matrixC0_0),
.matrixC0_1(matrixC0_1),
.matrixC0_2(matrixC0_2),
.matrixC0_3(matrixC0_3),
.matrixC0_4(matrixC0_4),
.matrixC0_5(matrixC0_5),
.matrixC0_6(matrixC0_6),
.matrixC0_7(matrixC0_7),
.matrixC0_8(matrixC0_8),
.matrixC0_9(matrixC0_9),
.matrixC0_10(matrixC0_10),
.matrixC0_11(matrixC0_11),
.matrixC0_12(matrixC0_12),
.matrixC0_13(matrixC0_13),
.matrixC0_14(matrixC0_14),
.matrixC0_15(matrixC0_15),
.matrixC0_16(matrixC0_16),
.matrixC0_17(matrixC0_17),
.matrixC0_18(matrixC0_18),
.matrixC0_19(matrixC0_19),
.matrixC0_20(matrixC0_20),
.matrixC0_21(matrixC0_21),
.matrixC0_22(matrixC0_22),
.matrixC0_23(matrixC0_23),
.matrixC0_24(matrixC0_24),
.matrixC0_25(matrixC0_25),
.matrixC0_26(matrixC0_26),
.matrixC0_27(matrixC0_27),
.matrixC0_28(matrixC0_28),
.matrixC0_29(matrixC0_29),
.matrixC0_30(matrixC0_30),
.matrixC0_31(matrixC0_31),
.matrixC1_0(matrixC1_0),
.matrixC1_1(matrixC1_1),
.matrixC1_2(matrixC1_2),
.matrixC1_3(matrixC1_3),
.matrixC1_4(matrixC1_4),
.matrixC1_5(matrixC1_5),
.matrixC1_6(matrixC1_6),
.matrixC1_7(matrixC1_7),
.matrixC1_8(matrixC1_8),
.matrixC1_9(matrixC1_9),
.matrixC1_10(matrixC1_10),
.matrixC1_11(matrixC1_11),
.matrixC1_12(matrixC1_12),
.matrixC1_13(matrixC1_13),
.matrixC1_14(matrixC1_14),
.matrixC1_15(matrixC1_15),
.matrixC1_16(matrixC1_16),
.matrixC1_17(matrixC1_17),
.matrixC1_18(matrixC1_18),
.matrixC1_19(matrixC1_19),
.matrixC1_20(matrixC1_20),
.matrixC1_21(matrixC1_21),
.matrixC1_22(matrixC1_22),
.matrixC1_23(matrixC1_23),
.matrixC1_24(matrixC1_24),
.matrixC1_25(matrixC1_25),
.matrixC1_26(matrixC1_26),
.matrixC1_27(matrixC1_27),
.matrixC1_28(matrixC1_28),
.matrixC1_29(matrixC1_29),
.matrixC1_30(matrixC1_30),
.matrixC1_31(matrixC1_31),
.matrixC2_0(matrixC2_0),
.matrixC2_1(matrixC2_1),
.matrixC2_2(matrixC2_2),
.matrixC2_3(matrixC2_3),
.matrixC2_4(matrixC2_4),
.matrixC2_5(matrixC2_5),
.matrixC2_6(matrixC2_6),
.matrixC2_7(matrixC2_7),
.matrixC2_8(matrixC2_8),
.matrixC2_9(matrixC2_9),
.matrixC2_10(matrixC2_10),
.matrixC2_11(matrixC2_11),
.matrixC2_12(matrixC2_12),
.matrixC2_13(matrixC2_13),
.matrixC2_14(matrixC2_14),
.matrixC2_15(matrixC2_15),
.matrixC2_16(matrixC2_16),
.matrixC2_17(matrixC2_17),
.matrixC2_18(matrixC2_18),
.matrixC2_19(matrixC2_19),
.matrixC2_20(matrixC2_20),
.matrixC2_21(matrixC2_21),
.matrixC2_22(matrixC2_22),
.matrixC2_23(matrixC2_23),
.matrixC2_24(matrixC2_24),
.matrixC2_25(matrixC2_25),
.matrixC2_26(matrixC2_26),
.matrixC2_27(matrixC2_27),
.matrixC2_28(matrixC2_28),
.matrixC2_29(matrixC2_29),
.matrixC2_30(matrixC2_30),
.matrixC2_31(matrixC2_31),
.matrixC3_0(matrixC3_0),
.matrixC3_1(matrixC3_1),
.matrixC3_2(matrixC3_2),
.matrixC3_3(matrixC3_3),
.matrixC3_4(matrixC3_4),
.matrixC3_5(matrixC3_5),
.matrixC3_6(matrixC3_6),
.matrixC3_7(matrixC3_7),
.matrixC3_8(matrixC3_8),
.matrixC3_9(matrixC3_9),
.matrixC3_10(matrixC3_10),
.matrixC3_11(matrixC3_11),
.matrixC3_12(matrixC3_12),
.matrixC3_13(matrixC3_13),
.matrixC3_14(matrixC3_14),
.matrixC3_15(matrixC3_15),
.matrixC3_16(matrixC3_16),
.matrixC3_17(matrixC3_17),
.matrixC3_18(matrixC3_18),
.matrixC3_19(matrixC3_19),
.matrixC3_20(matrixC3_20),
.matrixC3_21(matrixC3_21),
.matrixC3_22(matrixC3_22),
.matrixC3_23(matrixC3_23),
.matrixC3_24(matrixC3_24),
.matrixC3_25(matrixC3_25),
.matrixC3_26(matrixC3_26),
.matrixC3_27(matrixC3_27),
.matrixC3_28(matrixC3_28),
.matrixC3_29(matrixC3_29),
.matrixC3_30(matrixC3_30),
.matrixC3_31(matrixC3_31),
.matrixC4_0(matrixC4_0),
.matrixC4_1(matrixC4_1),
.matrixC4_2(matrixC4_2),
.matrixC4_3(matrixC4_3),
.matrixC4_4(matrixC4_4),
.matrixC4_5(matrixC4_5),
.matrixC4_6(matrixC4_6),
.matrixC4_7(matrixC4_7),
.matrixC4_8(matrixC4_8),
.matrixC4_9(matrixC4_9),
.matrixC4_10(matrixC4_10),
.matrixC4_11(matrixC4_11),
.matrixC4_12(matrixC4_12),
.matrixC4_13(matrixC4_13),
.matrixC4_14(matrixC4_14),
.matrixC4_15(matrixC4_15),
.matrixC4_16(matrixC4_16),
.matrixC4_17(matrixC4_17),
.matrixC4_18(matrixC4_18),
.matrixC4_19(matrixC4_19),
.matrixC4_20(matrixC4_20),
.matrixC4_21(matrixC4_21),
.matrixC4_22(matrixC4_22),
.matrixC4_23(matrixC4_23),
.matrixC4_24(matrixC4_24),
.matrixC4_25(matrixC4_25),
.matrixC4_26(matrixC4_26),
.matrixC4_27(matrixC4_27),
.matrixC4_28(matrixC4_28),
.matrixC4_29(matrixC4_29),
.matrixC4_30(matrixC4_30),
.matrixC4_31(matrixC4_31),
.matrixC5_0(matrixC5_0),
.matrixC5_1(matrixC5_1),
.matrixC5_2(matrixC5_2),
.matrixC5_3(matrixC5_3),
.matrixC5_4(matrixC5_4),
.matrixC5_5(matrixC5_5),
.matrixC5_6(matrixC5_6),
.matrixC5_7(matrixC5_7),
.matrixC5_8(matrixC5_8),
.matrixC5_9(matrixC5_9),
.matrixC5_10(matrixC5_10),
.matrixC5_11(matrixC5_11),
.matrixC5_12(matrixC5_12),
.matrixC5_13(matrixC5_13),
.matrixC5_14(matrixC5_14),
.matrixC5_15(matrixC5_15),
.matrixC5_16(matrixC5_16),
.matrixC5_17(matrixC5_17),
.matrixC5_18(matrixC5_18),
.matrixC5_19(matrixC5_19),
.matrixC5_20(matrixC5_20),
.matrixC5_21(matrixC5_21),
.matrixC5_22(matrixC5_22),
.matrixC5_23(matrixC5_23),
.matrixC5_24(matrixC5_24),
.matrixC5_25(matrixC5_25),
.matrixC5_26(matrixC5_26),
.matrixC5_27(matrixC5_27),
.matrixC5_28(matrixC5_28),
.matrixC5_29(matrixC5_29),
.matrixC5_30(matrixC5_30),
.matrixC5_31(matrixC5_31),
.matrixC6_0(matrixC6_0),
.matrixC6_1(matrixC6_1),
.matrixC6_2(matrixC6_2),
.matrixC6_3(matrixC6_3),
.matrixC6_4(matrixC6_4),
.matrixC6_5(matrixC6_5),
.matrixC6_6(matrixC6_6),
.matrixC6_7(matrixC6_7),
.matrixC6_8(matrixC6_8),
.matrixC6_9(matrixC6_9),
.matrixC6_10(matrixC6_10),
.matrixC6_11(matrixC6_11),
.matrixC6_12(matrixC6_12),
.matrixC6_13(matrixC6_13),
.matrixC6_14(matrixC6_14),
.matrixC6_15(matrixC6_15),
.matrixC6_16(matrixC6_16),
.matrixC6_17(matrixC6_17),
.matrixC6_18(matrixC6_18),
.matrixC6_19(matrixC6_19),
.matrixC6_20(matrixC6_20),
.matrixC6_21(matrixC6_21),
.matrixC6_22(matrixC6_22),
.matrixC6_23(matrixC6_23),
.matrixC6_24(matrixC6_24),
.matrixC6_25(matrixC6_25),
.matrixC6_26(matrixC6_26),
.matrixC6_27(matrixC6_27),
.matrixC6_28(matrixC6_28),
.matrixC6_29(matrixC6_29),
.matrixC6_30(matrixC6_30),
.matrixC6_31(matrixC6_31),
.matrixC7_0(matrixC7_0),
.matrixC7_1(matrixC7_1),
.matrixC7_2(matrixC7_2),
.matrixC7_3(matrixC7_3),
.matrixC7_4(matrixC7_4),
.matrixC7_5(matrixC7_5),
.matrixC7_6(matrixC7_6),
.matrixC7_7(matrixC7_7),
.matrixC7_8(matrixC7_8),
.matrixC7_9(matrixC7_9),
.matrixC7_10(matrixC7_10),
.matrixC7_11(matrixC7_11),
.matrixC7_12(matrixC7_12),
.matrixC7_13(matrixC7_13),
.matrixC7_14(matrixC7_14),
.matrixC7_15(matrixC7_15),
.matrixC7_16(matrixC7_16),
.matrixC7_17(matrixC7_17),
.matrixC7_18(matrixC7_18),
.matrixC7_19(matrixC7_19),
.matrixC7_20(matrixC7_20),
.matrixC7_21(matrixC7_21),
.matrixC7_22(matrixC7_22),
.matrixC7_23(matrixC7_23),
.matrixC7_24(matrixC7_24),
.matrixC7_25(matrixC7_25),
.matrixC7_26(matrixC7_26),
.matrixC7_27(matrixC7_27),
.matrixC7_28(matrixC7_28),
.matrixC7_29(matrixC7_29),
.matrixC7_30(matrixC7_30),
.matrixC7_31(matrixC7_31),
.matrixC8_0(matrixC8_0),
.matrixC8_1(matrixC8_1),
.matrixC8_2(matrixC8_2),
.matrixC8_3(matrixC8_3),
.matrixC8_4(matrixC8_4),
.matrixC8_5(matrixC8_5),
.matrixC8_6(matrixC8_6),
.matrixC8_7(matrixC8_7),
.matrixC8_8(matrixC8_8),
.matrixC8_9(matrixC8_9),
.matrixC8_10(matrixC8_10),
.matrixC8_11(matrixC8_11),
.matrixC8_12(matrixC8_12),
.matrixC8_13(matrixC8_13),
.matrixC8_14(matrixC8_14),
.matrixC8_15(matrixC8_15),
.matrixC8_16(matrixC8_16),
.matrixC8_17(matrixC8_17),
.matrixC8_18(matrixC8_18),
.matrixC8_19(matrixC8_19),
.matrixC8_20(matrixC8_20),
.matrixC8_21(matrixC8_21),
.matrixC8_22(matrixC8_22),
.matrixC8_23(matrixC8_23),
.matrixC8_24(matrixC8_24),
.matrixC8_25(matrixC8_25),
.matrixC8_26(matrixC8_26),
.matrixC8_27(matrixC8_27),
.matrixC8_28(matrixC8_28),
.matrixC8_29(matrixC8_29),
.matrixC8_30(matrixC8_30),
.matrixC8_31(matrixC8_31),
.matrixC9_0(matrixC9_0),
.matrixC9_1(matrixC9_1),
.matrixC9_2(matrixC9_2),
.matrixC9_3(matrixC9_3),
.matrixC9_4(matrixC9_4),
.matrixC9_5(matrixC9_5),
.matrixC9_6(matrixC9_6),
.matrixC9_7(matrixC9_7),
.matrixC9_8(matrixC9_8),
.matrixC9_9(matrixC9_9),
.matrixC9_10(matrixC9_10),
.matrixC9_11(matrixC9_11),
.matrixC9_12(matrixC9_12),
.matrixC9_13(matrixC9_13),
.matrixC9_14(matrixC9_14),
.matrixC9_15(matrixC9_15),
.matrixC9_16(matrixC9_16),
.matrixC9_17(matrixC9_17),
.matrixC9_18(matrixC9_18),
.matrixC9_19(matrixC9_19),
.matrixC9_20(matrixC9_20),
.matrixC9_21(matrixC9_21),
.matrixC9_22(matrixC9_22),
.matrixC9_23(matrixC9_23),
.matrixC9_24(matrixC9_24),
.matrixC9_25(matrixC9_25),
.matrixC9_26(matrixC9_26),
.matrixC9_27(matrixC9_27),
.matrixC9_28(matrixC9_28),
.matrixC9_29(matrixC9_29),
.matrixC9_30(matrixC9_30),
.matrixC9_31(matrixC9_31),
.matrixC10_0(matrixC10_0),
.matrixC10_1(matrixC10_1),
.matrixC10_2(matrixC10_2),
.matrixC10_3(matrixC10_3),
.matrixC10_4(matrixC10_4),
.matrixC10_5(matrixC10_5),
.matrixC10_6(matrixC10_6),
.matrixC10_7(matrixC10_7),
.matrixC10_8(matrixC10_8),
.matrixC10_9(matrixC10_9),
.matrixC10_10(matrixC10_10),
.matrixC10_11(matrixC10_11),
.matrixC10_12(matrixC10_12),
.matrixC10_13(matrixC10_13),
.matrixC10_14(matrixC10_14),
.matrixC10_15(matrixC10_15),
.matrixC10_16(matrixC10_16),
.matrixC10_17(matrixC10_17),
.matrixC10_18(matrixC10_18),
.matrixC10_19(matrixC10_19),
.matrixC10_20(matrixC10_20),
.matrixC10_21(matrixC10_21),
.matrixC10_22(matrixC10_22),
.matrixC10_23(matrixC10_23),
.matrixC10_24(matrixC10_24),
.matrixC10_25(matrixC10_25),
.matrixC10_26(matrixC10_26),
.matrixC10_27(matrixC10_27),
.matrixC10_28(matrixC10_28),
.matrixC10_29(matrixC10_29),
.matrixC10_30(matrixC10_30),
.matrixC10_31(matrixC10_31),
.matrixC11_0(matrixC11_0),
.matrixC11_1(matrixC11_1),
.matrixC11_2(matrixC11_2),
.matrixC11_3(matrixC11_3),
.matrixC11_4(matrixC11_4),
.matrixC11_5(matrixC11_5),
.matrixC11_6(matrixC11_6),
.matrixC11_7(matrixC11_7),
.matrixC11_8(matrixC11_8),
.matrixC11_9(matrixC11_9),
.matrixC11_10(matrixC11_10),
.matrixC11_11(matrixC11_11),
.matrixC11_12(matrixC11_12),
.matrixC11_13(matrixC11_13),
.matrixC11_14(matrixC11_14),
.matrixC11_15(matrixC11_15),
.matrixC11_16(matrixC11_16),
.matrixC11_17(matrixC11_17),
.matrixC11_18(matrixC11_18),
.matrixC11_19(matrixC11_19),
.matrixC11_20(matrixC11_20),
.matrixC11_21(matrixC11_21),
.matrixC11_22(matrixC11_22),
.matrixC11_23(matrixC11_23),
.matrixC11_24(matrixC11_24),
.matrixC11_25(matrixC11_25),
.matrixC11_26(matrixC11_26),
.matrixC11_27(matrixC11_27),
.matrixC11_28(matrixC11_28),
.matrixC11_29(matrixC11_29),
.matrixC11_30(matrixC11_30),
.matrixC11_31(matrixC11_31),
.matrixC12_0(matrixC12_0),
.matrixC12_1(matrixC12_1),
.matrixC12_2(matrixC12_2),
.matrixC12_3(matrixC12_3),
.matrixC12_4(matrixC12_4),
.matrixC12_5(matrixC12_5),
.matrixC12_6(matrixC12_6),
.matrixC12_7(matrixC12_7),
.matrixC12_8(matrixC12_8),
.matrixC12_9(matrixC12_9),
.matrixC12_10(matrixC12_10),
.matrixC12_11(matrixC12_11),
.matrixC12_12(matrixC12_12),
.matrixC12_13(matrixC12_13),
.matrixC12_14(matrixC12_14),
.matrixC12_15(matrixC12_15),
.matrixC12_16(matrixC12_16),
.matrixC12_17(matrixC12_17),
.matrixC12_18(matrixC12_18),
.matrixC12_19(matrixC12_19),
.matrixC12_20(matrixC12_20),
.matrixC12_21(matrixC12_21),
.matrixC12_22(matrixC12_22),
.matrixC12_23(matrixC12_23),
.matrixC12_24(matrixC12_24),
.matrixC12_25(matrixC12_25),
.matrixC12_26(matrixC12_26),
.matrixC12_27(matrixC12_27),
.matrixC12_28(matrixC12_28),
.matrixC12_29(matrixC12_29),
.matrixC12_30(matrixC12_30),
.matrixC12_31(matrixC12_31),
.matrixC13_0(matrixC13_0),
.matrixC13_1(matrixC13_1),
.matrixC13_2(matrixC13_2),
.matrixC13_3(matrixC13_3),
.matrixC13_4(matrixC13_4),
.matrixC13_5(matrixC13_5),
.matrixC13_6(matrixC13_6),
.matrixC13_7(matrixC13_7),
.matrixC13_8(matrixC13_8),
.matrixC13_9(matrixC13_9),
.matrixC13_10(matrixC13_10),
.matrixC13_11(matrixC13_11),
.matrixC13_12(matrixC13_12),
.matrixC13_13(matrixC13_13),
.matrixC13_14(matrixC13_14),
.matrixC13_15(matrixC13_15),
.matrixC13_16(matrixC13_16),
.matrixC13_17(matrixC13_17),
.matrixC13_18(matrixC13_18),
.matrixC13_19(matrixC13_19),
.matrixC13_20(matrixC13_20),
.matrixC13_21(matrixC13_21),
.matrixC13_22(matrixC13_22),
.matrixC13_23(matrixC13_23),
.matrixC13_24(matrixC13_24),
.matrixC13_25(matrixC13_25),
.matrixC13_26(matrixC13_26),
.matrixC13_27(matrixC13_27),
.matrixC13_28(matrixC13_28),
.matrixC13_29(matrixC13_29),
.matrixC13_30(matrixC13_30),
.matrixC13_31(matrixC13_31),
.matrixC14_0(matrixC14_0),
.matrixC14_1(matrixC14_1),
.matrixC14_2(matrixC14_2),
.matrixC14_3(matrixC14_3),
.matrixC14_4(matrixC14_4),
.matrixC14_5(matrixC14_5),
.matrixC14_6(matrixC14_6),
.matrixC14_7(matrixC14_7),
.matrixC14_8(matrixC14_8),
.matrixC14_9(matrixC14_9),
.matrixC14_10(matrixC14_10),
.matrixC14_11(matrixC14_11),
.matrixC14_12(matrixC14_12),
.matrixC14_13(matrixC14_13),
.matrixC14_14(matrixC14_14),
.matrixC14_15(matrixC14_15),
.matrixC14_16(matrixC14_16),
.matrixC14_17(matrixC14_17),
.matrixC14_18(matrixC14_18),
.matrixC14_19(matrixC14_19),
.matrixC14_20(matrixC14_20),
.matrixC14_21(matrixC14_21),
.matrixC14_22(matrixC14_22),
.matrixC14_23(matrixC14_23),
.matrixC14_24(matrixC14_24),
.matrixC14_25(matrixC14_25),
.matrixC14_26(matrixC14_26),
.matrixC14_27(matrixC14_27),
.matrixC14_28(matrixC14_28),
.matrixC14_29(matrixC14_29),
.matrixC14_30(matrixC14_30),
.matrixC14_31(matrixC14_31),
.matrixC15_0(matrixC15_0),
.matrixC15_1(matrixC15_1),
.matrixC15_2(matrixC15_2),
.matrixC15_3(matrixC15_3),
.matrixC15_4(matrixC15_4),
.matrixC15_5(matrixC15_5),
.matrixC15_6(matrixC15_6),
.matrixC15_7(matrixC15_7),
.matrixC15_8(matrixC15_8),
.matrixC15_9(matrixC15_9),
.matrixC15_10(matrixC15_10),
.matrixC15_11(matrixC15_11),
.matrixC15_12(matrixC15_12),
.matrixC15_13(matrixC15_13),
.matrixC15_14(matrixC15_14),
.matrixC15_15(matrixC15_15),
.matrixC15_16(matrixC15_16),
.matrixC15_17(matrixC15_17),
.matrixC15_18(matrixC15_18),
.matrixC15_19(matrixC15_19),
.matrixC15_20(matrixC15_20),
.matrixC15_21(matrixC15_21),
.matrixC15_22(matrixC15_22),
.matrixC15_23(matrixC15_23),
.matrixC15_24(matrixC15_24),
.matrixC15_25(matrixC15_25),
.matrixC15_26(matrixC15_26),
.matrixC15_27(matrixC15_27),
.matrixC15_28(matrixC15_28),
.matrixC15_29(matrixC15_29),
.matrixC15_30(matrixC15_30),
.matrixC15_31(matrixC15_31),
.matrixC16_0(matrixC16_0),
.matrixC16_1(matrixC16_1),
.matrixC16_2(matrixC16_2),
.matrixC16_3(matrixC16_3),
.matrixC16_4(matrixC16_4),
.matrixC16_5(matrixC16_5),
.matrixC16_6(matrixC16_6),
.matrixC16_7(matrixC16_7),
.matrixC16_8(matrixC16_8),
.matrixC16_9(matrixC16_9),
.matrixC16_10(matrixC16_10),
.matrixC16_11(matrixC16_11),
.matrixC16_12(matrixC16_12),
.matrixC16_13(matrixC16_13),
.matrixC16_14(matrixC16_14),
.matrixC16_15(matrixC16_15),
.matrixC16_16(matrixC16_16),
.matrixC16_17(matrixC16_17),
.matrixC16_18(matrixC16_18),
.matrixC16_19(matrixC16_19),
.matrixC16_20(matrixC16_20),
.matrixC16_21(matrixC16_21),
.matrixC16_22(matrixC16_22),
.matrixC16_23(matrixC16_23),
.matrixC16_24(matrixC16_24),
.matrixC16_25(matrixC16_25),
.matrixC16_26(matrixC16_26),
.matrixC16_27(matrixC16_27),
.matrixC16_28(matrixC16_28),
.matrixC16_29(matrixC16_29),
.matrixC16_30(matrixC16_30),
.matrixC16_31(matrixC16_31),
.matrixC17_0(matrixC17_0),
.matrixC17_1(matrixC17_1),
.matrixC17_2(matrixC17_2),
.matrixC17_3(matrixC17_3),
.matrixC17_4(matrixC17_4),
.matrixC17_5(matrixC17_5),
.matrixC17_6(matrixC17_6),
.matrixC17_7(matrixC17_7),
.matrixC17_8(matrixC17_8),
.matrixC17_9(matrixC17_9),
.matrixC17_10(matrixC17_10),
.matrixC17_11(matrixC17_11),
.matrixC17_12(matrixC17_12),
.matrixC17_13(matrixC17_13),
.matrixC17_14(matrixC17_14),
.matrixC17_15(matrixC17_15),
.matrixC17_16(matrixC17_16),
.matrixC17_17(matrixC17_17),
.matrixC17_18(matrixC17_18),
.matrixC17_19(matrixC17_19),
.matrixC17_20(matrixC17_20),
.matrixC17_21(matrixC17_21),
.matrixC17_22(matrixC17_22),
.matrixC17_23(matrixC17_23),
.matrixC17_24(matrixC17_24),
.matrixC17_25(matrixC17_25),
.matrixC17_26(matrixC17_26),
.matrixC17_27(matrixC17_27),
.matrixC17_28(matrixC17_28),
.matrixC17_29(matrixC17_29),
.matrixC17_30(matrixC17_30),
.matrixC17_31(matrixC17_31),
.matrixC18_0(matrixC18_0),
.matrixC18_1(matrixC18_1),
.matrixC18_2(matrixC18_2),
.matrixC18_3(matrixC18_3),
.matrixC18_4(matrixC18_4),
.matrixC18_5(matrixC18_5),
.matrixC18_6(matrixC18_6),
.matrixC18_7(matrixC18_7),
.matrixC18_8(matrixC18_8),
.matrixC18_9(matrixC18_9),
.matrixC18_10(matrixC18_10),
.matrixC18_11(matrixC18_11),
.matrixC18_12(matrixC18_12),
.matrixC18_13(matrixC18_13),
.matrixC18_14(matrixC18_14),
.matrixC18_15(matrixC18_15),
.matrixC18_16(matrixC18_16),
.matrixC18_17(matrixC18_17),
.matrixC18_18(matrixC18_18),
.matrixC18_19(matrixC18_19),
.matrixC18_20(matrixC18_20),
.matrixC18_21(matrixC18_21),
.matrixC18_22(matrixC18_22),
.matrixC18_23(matrixC18_23),
.matrixC18_24(matrixC18_24),
.matrixC18_25(matrixC18_25),
.matrixC18_26(matrixC18_26),
.matrixC18_27(matrixC18_27),
.matrixC18_28(matrixC18_28),
.matrixC18_29(matrixC18_29),
.matrixC18_30(matrixC18_30),
.matrixC18_31(matrixC18_31),
.matrixC19_0(matrixC19_0),
.matrixC19_1(matrixC19_1),
.matrixC19_2(matrixC19_2),
.matrixC19_3(matrixC19_3),
.matrixC19_4(matrixC19_4),
.matrixC19_5(matrixC19_5),
.matrixC19_6(matrixC19_6),
.matrixC19_7(matrixC19_7),
.matrixC19_8(matrixC19_8),
.matrixC19_9(matrixC19_9),
.matrixC19_10(matrixC19_10),
.matrixC19_11(matrixC19_11),
.matrixC19_12(matrixC19_12),
.matrixC19_13(matrixC19_13),
.matrixC19_14(matrixC19_14),
.matrixC19_15(matrixC19_15),
.matrixC19_16(matrixC19_16),
.matrixC19_17(matrixC19_17),
.matrixC19_18(matrixC19_18),
.matrixC19_19(matrixC19_19),
.matrixC19_20(matrixC19_20),
.matrixC19_21(matrixC19_21),
.matrixC19_22(matrixC19_22),
.matrixC19_23(matrixC19_23),
.matrixC19_24(matrixC19_24),
.matrixC19_25(matrixC19_25),
.matrixC19_26(matrixC19_26),
.matrixC19_27(matrixC19_27),
.matrixC19_28(matrixC19_28),
.matrixC19_29(matrixC19_29),
.matrixC19_30(matrixC19_30),
.matrixC19_31(matrixC19_31),
.matrixC20_0(matrixC20_0),
.matrixC20_1(matrixC20_1),
.matrixC20_2(matrixC20_2),
.matrixC20_3(matrixC20_3),
.matrixC20_4(matrixC20_4),
.matrixC20_5(matrixC20_5),
.matrixC20_6(matrixC20_6),
.matrixC20_7(matrixC20_7),
.matrixC20_8(matrixC20_8),
.matrixC20_9(matrixC20_9),
.matrixC20_10(matrixC20_10),
.matrixC20_11(matrixC20_11),
.matrixC20_12(matrixC20_12),
.matrixC20_13(matrixC20_13),
.matrixC20_14(matrixC20_14),
.matrixC20_15(matrixC20_15),
.matrixC20_16(matrixC20_16),
.matrixC20_17(matrixC20_17),
.matrixC20_18(matrixC20_18),
.matrixC20_19(matrixC20_19),
.matrixC20_20(matrixC20_20),
.matrixC20_21(matrixC20_21),
.matrixC20_22(matrixC20_22),
.matrixC20_23(matrixC20_23),
.matrixC20_24(matrixC20_24),
.matrixC20_25(matrixC20_25),
.matrixC20_26(matrixC20_26),
.matrixC20_27(matrixC20_27),
.matrixC20_28(matrixC20_28),
.matrixC20_29(matrixC20_29),
.matrixC20_30(matrixC20_30),
.matrixC20_31(matrixC20_31),
.matrixC21_0(matrixC21_0),
.matrixC21_1(matrixC21_1),
.matrixC21_2(matrixC21_2),
.matrixC21_3(matrixC21_3),
.matrixC21_4(matrixC21_4),
.matrixC21_5(matrixC21_5),
.matrixC21_6(matrixC21_6),
.matrixC21_7(matrixC21_7),
.matrixC21_8(matrixC21_8),
.matrixC21_9(matrixC21_9),
.matrixC21_10(matrixC21_10),
.matrixC21_11(matrixC21_11),
.matrixC21_12(matrixC21_12),
.matrixC21_13(matrixC21_13),
.matrixC21_14(matrixC21_14),
.matrixC21_15(matrixC21_15),
.matrixC21_16(matrixC21_16),
.matrixC21_17(matrixC21_17),
.matrixC21_18(matrixC21_18),
.matrixC21_19(matrixC21_19),
.matrixC21_20(matrixC21_20),
.matrixC21_21(matrixC21_21),
.matrixC21_22(matrixC21_22),
.matrixC21_23(matrixC21_23),
.matrixC21_24(matrixC21_24),
.matrixC21_25(matrixC21_25),
.matrixC21_26(matrixC21_26),
.matrixC21_27(matrixC21_27),
.matrixC21_28(matrixC21_28),
.matrixC21_29(matrixC21_29),
.matrixC21_30(matrixC21_30),
.matrixC21_31(matrixC21_31),
.matrixC22_0(matrixC22_0),
.matrixC22_1(matrixC22_1),
.matrixC22_2(matrixC22_2),
.matrixC22_3(matrixC22_3),
.matrixC22_4(matrixC22_4),
.matrixC22_5(matrixC22_5),
.matrixC22_6(matrixC22_6),
.matrixC22_7(matrixC22_7),
.matrixC22_8(matrixC22_8),
.matrixC22_9(matrixC22_9),
.matrixC22_10(matrixC22_10),
.matrixC22_11(matrixC22_11),
.matrixC22_12(matrixC22_12),
.matrixC22_13(matrixC22_13),
.matrixC22_14(matrixC22_14),
.matrixC22_15(matrixC22_15),
.matrixC22_16(matrixC22_16),
.matrixC22_17(matrixC22_17),
.matrixC22_18(matrixC22_18),
.matrixC22_19(matrixC22_19),
.matrixC22_20(matrixC22_20),
.matrixC22_21(matrixC22_21),
.matrixC22_22(matrixC22_22),
.matrixC22_23(matrixC22_23),
.matrixC22_24(matrixC22_24),
.matrixC22_25(matrixC22_25),
.matrixC22_26(matrixC22_26),
.matrixC22_27(matrixC22_27),
.matrixC22_28(matrixC22_28),
.matrixC22_29(matrixC22_29),
.matrixC22_30(matrixC22_30),
.matrixC22_31(matrixC22_31),
.matrixC23_0(matrixC23_0),
.matrixC23_1(matrixC23_1),
.matrixC23_2(matrixC23_2),
.matrixC23_3(matrixC23_3),
.matrixC23_4(matrixC23_4),
.matrixC23_5(matrixC23_5),
.matrixC23_6(matrixC23_6),
.matrixC23_7(matrixC23_7),
.matrixC23_8(matrixC23_8),
.matrixC23_9(matrixC23_9),
.matrixC23_10(matrixC23_10),
.matrixC23_11(matrixC23_11),
.matrixC23_12(matrixC23_12),
.matrixC23_13(matrixC23_13),
.matrixC23_14(matrixC23_14),
.matrixC23_15(matrixC23_15),
.matrixC23_16(matrixC23_16),
.matrixC23_17(matrixC23_17),
.matrixC23_18(matrixC23_18),
.matrixC23_19(matrixC23_19),
.matrixC23_20(matrixC23_20),
.matrixC23_21(matrixC23_21),
.matrixC23_22(matrixC23_22),
.matrixC23_23(matrixC23_23),
.matrixC23_24(matrixC23_24),
.matrixC23_25(matrixC23_25),
.matrixC23_26(matrixC23_26),
.matrixC23_27(matrixC23_27),
.matrixC23_28(matrixC23_28),
.matrixC23_29(matrixC23_29),
.matrixC23_30(matrixC23_30),
.matrixC23_31(matrixC23_31),
.matrixC24_0(matrixC24_0),
.matrixC24_1(matrixC24_1),
.matrixC24_2(matrixC24_2),
.matrixC24_3(matrixC24_3),
.matrixC24_4(matrixC24_4),
.matrixC24_5(matrixC24_5),
.matrixC24_6(matrixC24_6),
.matrixC24_7(matrixC24_7),
.matrixC24_8(matrixC24_8),
.matrixC24_9(matrixC24_9),
.matrixC24_10(matrixC24_10),
.matrixC24_11(matrixC24_11),
.matrixC24_12(matrixC24_12),
.matrixC24_13(matrixC24_13),
.matrixC24_14(matrixC24_14),
.matrixC24_15(matrixC24_15),
.matrixC24_16(matrixC24_16),
.matrixC24_17(matrixC24_17),
.matrixC24_18(matrixC24_18),
.matrixC24_19(matrixC24_19),
.matrixC24_20(matrixC24_20),
.matrixC24_21(matrixC24_21),
.matrixC24_22(matrixC24_22),
.matrixC24_23(matrixC24_23),
.matrixC24_24(matrixC24_24),
.matrixC24_25(matrixC24_25),
.matrixC24_26(matrixC24_26),
.matrixC24_27(matrixC24_27),
.matrixC24_28(matrixC24_28),
.matrixC24_29(matrixC24_29),
.matrixC24_30(matrixC24_30),
.matrixC24_31(matrixC24_31),
.matrixC25_0(matrixC25_0),
.matrixC25_1(matrixC25_1),
.matrixC25_2(matrixC25_2),
.matrixC25_3(matrixC25_3),
.matrixC25_4(matrixC25_4),
.matrixC25_5(matrixC25_5),
.matrixC25_6(matrixC25_6),
.matrixC25_7(matrixC25_7),
.matrixC25_8(matrixC25_8),
.matrixC25_9(matrixC25_9),
.matrixC25_10(matrixC25_10),
.matrixC25_11(matrixC25_11),
.matrixC25_12(matrixC25_12),
.matrixC25_13(matrixC25_13),
.matrixC25_14(matrixC25_14),
.matrixC25_15(matrixC25_15),
.matrixC25_16(matrixC25_16),
.matrixC25_17(matrixC25_17),
.matrixC25_18(matrixC25_18),
.matrixC25_19(matrixC25_19),
.matrixC25_20(matrixC25_20),
.matrixC25_21(matrixC25_21),
.matrixC25_22(matrixC25_22),
.matrixC25_23(matrixC25_23),
.matrixC25_24(matrixC25_24),
.matrixC25_25(matrixC25_25),
.matrixC25_26(matrixC25_26),
.matrixC25_27(matrixC25_27),
.matrixC25_28(matrixC25_28),
.matrixC25_29(matrixC25_29),
.matrixC25_30(matrixC25_30),
.matrixC25_31(matrixC25_31),
.matrixC26_0(matrixC26_0),
.matrixC26_1(matrixC26_1),
.matrixC26_2(matrixC26_2),
.matrixC26_3(matrixC26_3),
.matrixC26_4(matrixC26_4),
.matrixC26_5(matrixC26_5),
.matrixC26_6(matrixC26_6),
.matrixC26_7(matrixC26_7),
.matrixC26_8(matrixC26_8),
.matrixC26_9(matrixC26_9),
.matrixC26_10(matrixC26_10),
.matrixC26_11(matrixC26_11),
.matrixC26_12(matrixC26_12),
.matrixC26_13(matrixC26_13),
.matrixC26_14(matrixC26_14),
.matrixC26_15(matrixC26_15),
.matrixC26_16(matrixC26_16),
.matrixC26_17(matrixC26_17),
.matrixC26_18(matrixC26_18),
.matrixC26_19(matrixC26_19),
.matrixC26_20(matrixC26_20),
.matrixC26_21(matrixC26_21),
.matrixC26_22(matrixC26_22),
.matrixC26_23(matrixC26_23),
.matrixC26_24(matrixC26_24),
.matrixC26_25(matrixC26_25),
.matrixC26_26(matrixC26_26),
.matrixC26_27(matrixC26_27),
.matrixC26_28(matrixC26_28),
.matrixC26_29(matrixC26_29),
.matrixC26_30(matrixC26_30),
.matrixC26_31(matrixC26_31),
.matrixC27_0(matrixC27_0),
.matrixC27_1(matrixC27_1),
.matrixC27_2(matrixC27_2),
.matrixC27_3(matrixC27_3),
.matrixC27_4(matrixC27_4),
.matrixC27_5(matrixC27_5),
.matrixC27_6(matrixC27_6),
.matrixC27_7(matrixC27_7),
.matrixC27_8(matrixC27_8),
.matrixC27_9(matrixC27_9),
.matrixC27_10(matrixC27_10),
.matrixC27_11(matrixC27_11),
.matrixC27_12(matrixC27_12),
.matrixC27_13(matrixC27_13),
.matrixC27_14(matrixC27_14),
.matrixC27_15(matrixC27_15),
.matrixC27_16(matrixC27_16),
.matrixC27_17(matrixC27_17),
.matrixC27_18(matrixC27_18),
.matrixC27_19(matrixC27_19),
.matrixC27_20(matrixC27_20),
.matrixC27_21(matrixC27_21),
.matrixC27_22(matrixC27_22),
.matrixC27_23(matrixC27_23),
.matrixC27_24(matrixC27_24),
.matrixC27_25(matrixC27_25),
.matrixC27_26(matrixC27_26),
.matrixC27_27(matrixC27_27),
.matrixC27_28(matrixC27_28),
.matrixC27_29(matrixC27_29),
.matrixC27_30(matrixC27_30),
.matrixC27_31(matrixC27_31),
.matrixC28_0(matrixC28_0),
.matrixC28_1(matrixC28_1),
.matrixC28_2(matrixC28_2),
.matrixC28_3(matrixC28_3),
.matrixC28_4(matrixC28_4),
.matrixC28_5(matrixC28_5),
.matrixC28_6(matrixC28_6),
.matrixC28_7(matrixC28_7),
.matrixC28_8(matrixC28_8),
.matrixC28_9(matrixC28_9),
.matrixC28_10(matrixC28_10),
.matrixC28_11(matrixC28_11),
.matrixC28_12(matrixC28_12),
.matrixC28_13(matrixC28_13),
.matrixC28_14(matrixC28_14),
.matrixC28_15(matrixC28_15),
.matrixC28_16(matrixC28_16),
.matrixC28_17(matrixC28_17),
.matrixC28_18(matrixC28_18),
.matrixC28_19(matrixC28_19),
.matrixC28_20(matrixC28_20),
.matrixC28_21(matrixC28_21),
.matrixC28_22(matrixC28_22),
.matrixC28_23(matrixC28_23),
.matrixC28_24(matrixC28_24),
.matrixC28_25(matrixC28_25),
.matrixC28_26(matrixC28_26),
.matrixC28_27(matrixC28_27),
.matrixC28_28(matrixC28_28),
.matrixC28_29(matrixC28_29),
.matrixC28_30(matrixC28_30),
.matrixC28_31(matrixC28_31),
.matrixC29_0(matrixC29_0),
.matrixC29_1(matrixC29_1),
.matrixC29_2(matrixC29_2),
.matrixC29_3(matrixC29_3),
.matrixC29_4(matrixC29_4),
.matrixC29_5(matrixC29_5),
.matrixC29_6(matrixC29_6),
.matrixC29_7(matrixC29_7),
.matrixC29_8(matrixC29_8),
.matrixC29_9(matrixC29_9),
.matrixC29_10(matrixC29_10),
.matrixC29_11(matrixC29_11),
.matrixC29_12(matrixC29_12),
.matrixC29_13(matrixC29_13),
.matrixC29_14(matrixC29_14),
.matrixC29_15(matrixC29_15),
.matrixC29_16(matrixC29_16),
.matrixC29_17(matrixC29_17),
.matrixC29_18(matrixC29_18),
.matrixC29_19(matrixC29_19),
.matrixC29_20(matrixC29_20),
.matrixC29_21(matrixC29_21),
.matrixC29_22(matrixC29_22),
.matrixC29_23(matrixC29_23),
.matrixC29_24(matrixC29_24),
.matrixC29_25(matrixC29_25),
.matrixC29_26(matrixC29_26),
.matrixC29_27(matrixC29_27),
.matrixC29_28(matrixC29_28),
.matrixC29_29(matrixC29_29),
.matrixC29_30(matrixC29_30),
.matrixC29_31(matrixC29_31),
.matrixC30_0(matrixC30_0),
.matrixC30_1(matrixC30_1),
.matrixC30_2(matrixC30_2),
.matrixC30_3(matrixC30_3),
.matrixC30_4(matrixC30_4),
.matrixC30_5(matrixC30_5),
.matrixC30_6(matrixC30_6),
.matrixC30_7(matrixC30_7),
.matrixC30_8(matrixC30_8),
.matrixC30_9(matrixC30_9),
.matrixC30_10(matrixC30_10),
.matrixC30_11(matrixC30_11),
.matrixC30_12(matrixC30_12),
.matrixC30_13(matrixC30_13),
.matrixC30_14(matrixC30_14),
.matrixC30_15(matrixC30_15),
.matrixC30_16(matrixC30_16),
.matrixC30_17(matrixC30_17),
.matrixC30_18(matrixC30_18),
.matrixC30_19(matrixC30_19),
.matrixC30_20(matrixC30_20),
.matrixC30_21(matrixC30_21),
.matrixC30_22(matrixC30_22),
.matrixC30_23(matrixC30_23),
.matrixC30_24(matrixC30_24),
.matrixC30_25(matrixC30_25),
.matrixC30_26(matrixC30_26),
.matrixC30_27(matrixC30_27),
.matrixC30_28(matrixC30_28),
.matrixC30_29(matrixC30_29),
.matrixC30_30(matrixC30_30),
.matrixC30_31(matrixC30_31),
.matrixC31_0(matrixC31_0),
.matrixC31_1(matrixC31_1),
.matrixC31_2(matrixC31_2),
.matrixC31_3(matrixC31_3),
.matrixC31_4(matrixC31_4),
.matrixC31_5(matrixC31_5),
.matrixC31_6(matrixC31_6),
.matrixC31_7(matrixC31_7),
.matrixC31_8(matrixC31_8),
.matrixC31_9(matrixC31_9),
.matrixC31_10(matrixC31_10),
.matrixC31_11(matrixC31_11),
.matrixC31_12(matrixC31_12),
.matrixC31_13(matrixC31_13),
.matrixC31_14(matrixC31_14),
.matrixC31_15(matrixC31_15),
.matrixC31_16(matrixC31_16),
.matrixC31_17(matrixC31_17),
.matrixC31_18(matrixC31_18),
.matrixC31_19(matrixC31_19),
.matrixC31_20(matrixC31_20),
.matrixC31_21(matrixC31_21),
.matrixC31_22(matrixC31_22),
.matrixC31_23(matrixC31_23),
.matrixC31_24(matrixC31_24),
.matrixC31_25(matrixC31_25),
.matrixC31_26(matrixC31_26),
.matrixC31_27(matrixC31_27),
.matrixC31_28(matrixC31_28),
.matrixC31_29(matrixC31_29),
.matrixC31_30(matrixC31_30),
.matrixC31_31(matrixC31_31),

.a_data_out(a_data_out),
.b_data_out(b_data_out)
);

endmodule


//////////////////////////////////////////////////////////////////////////
// Output logic
//////////////////////////////////////////////////////////////////////////
module output_logic(
start_mat_mul,
done_mat_mul,
address_mat_c,
address_stride_c,
c_data_in,
c_data_out, //Data values going out to next matmul - systolic shifting
c_addr,
c_data_available,
clk_cnt,
row_latch_en,

final_mat_mul_size,
  matrixC0_0,
matrixC0_1,
matrixC0_2,
matrixC0_3,
matrixC0_4,
matrixC0_5,
matrixC0_6,
matrixC0_7,
matrixC0_8,
matrixC0_9,
matrixC0_10,
matrixC0_11,
matrixC0_12,
matrixC0_13,
matrixC0_14,
matrixC0_15,
matrixC0_16,
matrixC0_17,
matrixC0_18,
matrixC0_19,
matrixC0_20,
matrixC0_21,
matrixC0_22,
matrixC0_23,
matrixC0_24,
matrixC0_25,
matrixC0_26,
matrixC0_27,
matrixC0_28,
matrixC0_29,
matrixC0_30,
matrixC0_31,
matrixC1_0,
matrixC1_1,
matrixC1_2,
matrixC1_3,
matrixC1_4,
matrixC1_5,
matrixC1_6,
matrixC1_7,
matrixC1_8,
matrixC1_9,
matrixC1_10,
matrixC1_11,
matrixC1_12,
matrixC1_13,
matrixC1_14,
matrixC1_15,
matrixC1_16,
matrixC1_17,
matrixC1_18,
matrixC1_19,
matrixC1_20,
matrixC1_21,
matrixC1_22,
matrixC1_23,
matrixC1_24,
matrixC1_25,
matrixC1_26,
matrixC1_27,
matrixC1_28,
matrixC1_29,
matrixC1_30,
matrixC1_31,
matrixC2_0,
matrixC2_1,
matrixC2_2,
matrixC2_3,
matrixC2_4,
matrixC2_5,
matrixC2_6,
matrixC2_7,
matrixC2_8,
matrixC2_9,
matrixC2_10,
matrixC2_11,
matrixC2_12,
matrixC2_13,
matrixC2_14,
matrixC2_15,
matrixC2_16,
matrixC2_17,
matrixC2_18,
matrixC2_19,
matrixC2_20,
matrixC2_21,
matrixC2_22,
matrixC2_23,
matrixC2_24,
matrixC2_25,
matrixC2_26,
matrixC2_27,
matrixC2_28,
matrixC2_29,
matrixC2_30,
matrixC2_31,
matrixC3_0,
matrixC3_1,
matrixC3_2,
matrixC3_3,
matrixC3_4,
matrixC3_5,
matrixC3_6,
matrixC3_7,
matrixC3_8,
matrixC3_9,
matrixC3_10,
matrixC3_11,
matrixC3_12,
matrixC3_13,
matrixC3_14,
matrixC3_15,
matrixC3_16,
matrixC3_17,
matrixC3_18,
matrixC3_19,
matrixC3_20,
matrixC3_21,
matrixC3_22,
matrixC3_23,
matrixC3_24,
matrixC3_25,
matrixC3_26,
matrixC3_27,
matrixC3_28,
matrixC3_29,
matrixC3_30,
matrixC3_31,
matrixC4_0,
matrixC4_1,
matrixC4_2,
matrixC4_3,
matrixC4_4,
matrixC4_5,
matrixC4_6,
matrixC4_7,
matrixC4_8,
matrixC4_9,
matrixC4_10,
matrixC4_11,
matrixC4_12,
matrixC4_13,
matrixC4_14,
matrixC4_15,
matrixC4_16,
matrixC4_17,
matrixC4_18,
matrixC4_19,
matrixC4_20,
matrixC4_21,
matrixC4_22,
matrixC4_23,
matrixC4_24,
matrixC4_25,
matrixC4_26,
matrixC4_27,
matrixC4_28,
matrixC4_29,
matrixC4_30,
matrixC4_31,
matrixC5_0,
matrixC5_1,
matrixC5_2,
matrixC5_3,
matrixC5_4,
matrixC5_5,
matrixC5_6,
matrixC5_7,
matrixC5_8,
matrixC5_9,
matrixC5_10,
matrixC5_11,
matrixC5_12,
matrixC5_13,
matrixC5_14,
matrixC5_15,
matrixC5_16,
matrixC5_17,
matrixC5_18,
matrixC5_19,
matrixC5_20,
matrixC5_21,
matrixC5_22,
matrixC5_23,
matrixC5_24,
matrixC5_25,
matrixC5_26,
matrixC5_27,
matrixC5_28,
matrixC5_29,
matrixC5_30,
matrixC5_31,
matrixC6_0,
matrixC6_1,
matrixC6_2,
matrixC6_3,
matrixC6_4,
matrixC6_5,
matrixC6_6,
matrixC6_7,
matrixC6_8,
matrixC6_9,
matrixC6_10,
matrixC6_11,
matrixC6_12,
matrixC6_13,
matrixC6_14,
matrixC6_15,
matrixC6_16,
matrixC6_17,
matrixC6_18,
matrixC6_19,
matrixC6_20,
matrixC6_21,
matrixC6_22,
matrixC6_23,
matrixC6_24,
matrixC6_25,
matrixC6_26,
matrixC6_27,
matrixC6_28,
matrixC6_29,
matrixC6_30,
matrixC6_31,
matrixC7_0,
matrixC7_1,
matrixC7_2,
matrixC7_3,
matrixC7_4,
matrixC7_5,
matrixC7_6,
matrixC7_7,
matrixC7_8,
matrixC7_9,
matrixC7_10,
matrixC7_11,
matrixC7_12,
matrixC7_13,
matrixC7_14,
matrixC7_15,
matrixC7_16,
matrixC7_17,
matrixC7_18,
matrixC7_19,
matrixC7_20,
matrixC7_21,
matrixC7_22,
matrixC7_23,
matrixC7_24,
matrixC7_25,
matrixC7_26,
matrixC7_27,
matrixC7_28,
matrixC7_29,
matrixC7_30,
matrixC7_31,
matrixC8_0,
matrixC8_1,
matrixC8_2,
matrixC8_3,
matrixC8_4,
matrixC8_5,
matrixC8_6,
matrixC8_7,
matrixC8_8,
matrixC8_9,
matrixC8_10,
matrixC8_11,
matrixC8_12,
matrixC8_13,
matrixC8_14,
matrixC8_15,
matrixC8_16,
matrixC8_17,
matrixC8_18,
matrixC8_19,
matrixC8_20,
matrixC8_21,
matrixC8_22,
matrixC8_23,
matrixC8_24,
matrixC8_25,
matrixC8_26,
matrixC8_27,
matrixC8_28,
matrixC8_29,
matrixC8_30,
matrixC8_31,
matrixC9_0,
matrixC9_1,
matrixC9_2,
matrixC9_3,
matrixC9_4,
matrixC9_5,
matrixC9_6,
matrixC9_7,
matrixC9_8,
matrixC9_9,
matrixC9_10,
matrixC9_11,
matrixC9_12,
matrixC9_13,
matrixC9_14,
matrixC9_15,
matrixC9_16,
matrixC9_17,
matrixC9_18,
matrixC9_19,
matrixC9_20,
matrixC9_21,
matrixC9_22,
matrixC9_23,
matrixC9_24,
matrixC9_25,
matrixC9_26,
matrixC9_27,
matrixC9_28,
matrixC9_29,
matrixC9_30,
matrixC9_31,
matrixC10_0,
matrixC10_1,
matrixC10_2,
matrixC10_3,
matrixC10_4,
matrixC10_5,
matrixC10_6,
matrixC10_7,
matrixC10_8,
matrixC10_9,
matrixC10_10,
matrixC10_11,
matrixC10_12,
matrixC10_13,
matrixC10_14,
matrixC10_15,
matrixC10_16,
matrixC10_17,
matrixC10_18,
matrixC10_19,
matrixC10_20,
matrixC10_21,
matrixC10_22,
matrixC10_23,
matrixC10_24,
matrixC10_25,
matrixC10_26,
matrixC10_27,
matrixC10_28,
matrixC10_29,
matrixC10_30,
matrixC10_31,
matrixC11_0,
matrixC11_1,
matrixC11_2,
matrixC11_3,
matrixC11_4,
matrixC11_5,
matrixC11_6,
matrixC11_7,
matrixC11_8,
matrixC11_9,
matrixC11_10,
matrixC11_11,
matrixC11_12,
matrixC11_13,
matrixC11_14,
matrixC11_15,
matrixC11_16,
matrixC11_17,
matrixC11_18,
matrixC11_19,
matrixC11_20,
matrixC11_21,
matrixC11_22,
matrixC11_23,
matrixC11_24,
matrixC11_25,
matrixC11_26,
matrixC11_27,
matrixC11_28,
matrixC11_29,
matrixC11_30,
matrixC11_31,
matrixC12_0,
matrixC12_1,
matrixC12_2,
matrixC12_3,
matrixC12_4,
matrixC12_5,
matrixC12_6,
matrixC12_7,
matrixC12_8,
matrixC12_9,
matrixC12_10,
matrixC12_11,
matrixC12_12,
matrixC12_13,
matrixC12_14,
matrixC12_15,
matrixC12_16,
matrixC12_17,
matrixC12_18,
matrixC12_19,
matrixC12_20,
matrixC12_21,
matrixC12_22,
matrixC12_23,
matrixC12_24,
matrixC12_25,
matrixC12_26,
matrixC12_27,
matrixC12_28,
matrixC12_29,
matrixC12_30,
matrixC12_31,
matrixC13_0,
matrixC13_1,
matrixC13_2,
matrixC13_3,
matrixC13_4,
matrixC13_5,
matrixC13_6,
matrixC13_7,
matrixC13_8,
matrixC13_9,
matrixC13_10,
matrixC13_11,
matrixC13_12,
matrixC13_13,
matrixC13_14,
matrixC13_15,
matrixC13_16,
matrixC13_17,
matrixC13_18,
matrixC13_19,
matrixC13_20,
matrixC13_21,
matrixC13_22,
matrixC13_23,
matrixC13_24,
matrixC13_25,
matrixC13_26,
matrixC13_27,
matrixC13_28,
matrixC13_29,
matrixC13_30,
matrixC13_31,
matrixC14_0,
matrixC14_1,
matrixC14_2,
matrixC14_3,
matrixC14_4,
matrixC14_5,
matrixC14_6,
matrixC14_7,
matrixC14_8,
matrixC14_9,
matrixC14_10,
matrixC14_11,
matrixC14_12,
matrixC14_13,
matrixC14_14,
matrixC14_15,
matrixC14_16,
matrixC14_17,
matrixC14_18,
matrixC14_19,
matrixC14_20,
matrixC14_21,
matrixC14_22,
matrixC14_23,
matrixC14_24,
matrixC14_25,
matrixC14_26,
matrixC14_27,
matrixC14_28,
matrixC14_29,
matrixC14_30,
matrixC14_31,
matrixC15_0,
matrixC15_1,
matrixC15_2,
matrixC15_3,
matrixC15_4,
matrixC15_5,
matrixC15_6,
matrixC15_7,
matrixC15_8,
matrixC15_9,
matrixC15_10,
matrixC15_11,
matrixC15_12,
matrixC15_13,
matrixC15_14,
matrixC15_15,
matrixC15_16,
matrixC15_17,
matrixC15_18,
matrixC15_19,
matrixC15_20,
matrixC15_21,
matrixC15_22,
matrixC15_23,
matrixC15_24,
matrixC15_25,
matrixC15_26,
matrixC15_27,
matrixC15_28,
matrixC15_29,
matrixC15_30,
matrixC15_31,
matrixC16_0,
matrixC16_1,
matrixC16_2,
matrixC16_3,
matrixC16_4,
matrixC16_5,
matrixC16_6,
matrixC16_7,
matrixC16_8,
matrixC16_9,
matrixC16_10,
matrixC16_11,
matrixC16_12,
matrixC16_13,
matrixC16_14,
matrixC16_15,
matrixC16_16,
matrixC16_17,
matrixC16_18,
matrixC16_19,
matrixC16_20,
matrixC16_21,
matrixC16_22,
matrixC16_23,
matrixC16_24,
matrixC16_25,
matrixC16_26,
matrixC16_27,
matrixC16_28,
matrixC16_29,
matrixC16_30,
matrixC16_31,
matrixC17_0,
matrixC17_1,
matrixC17_2,
matrixC17_3,
matrixC17_4,
matrixC17_5,
matrixC17_6,
matrixC17_7,
matrixC17_8,
matrixC17_9,
matrixC17_10,
matrixC17_11,
matrixC17_12,
matrixC17_13,
matrixC17_14,
matrixC17_15,
matrixC17_16,
matrixC17_17,
matrixC17_18,
matrixC17_19,
matrixC17_20,
matrixC17_21,
matrixC17_22,
matrixC17_23,
matrixC17_24,
matrixC17_25,
matrixC17_26,
matrixC17_27,
matrixC17_28,
matrixC17_29,
matrixC17_30,
matrixC17_31,
matrixC18_0,
matrixC18_1,
matrixC18_2,
matrixC18_3,
matrixC18_4,
matrixC18_5,
matrixC18_6,
matrixC18_7,
matrixC18_8,
matrixC18_9,
matrixC18_10,
matrixC18_11,
matrixC18_12,
matrixC18_13,
matrixC18_14,
matrixC18_15,
matrixC18_16,
matrixC18_17,
matrixC18_18,
matrixC18_19,
matrixC18_20,
matrixC18_21,
matrixC18_22,
matrixC18_23,
matrixC18_24,
matrixC18_25,
matrixC18_26,
matrixC18_27,
matrixC18_28,
matrixC18_29,
matrixC18_30,
matrixC18_31,
matrixC19_0,
matrixC19_1,
matrixC19_2,
matrixC19_3,
matrixC19_4,
matrixC19_5,
matrixC19_6,
matrixC19_7,
matrixC19_8,
matrixC19_9,
matrixC19_10,
matrixC19_11,
matrixC19_12,
matrixC19_13,
matrixC19_14,
matrixC19_15,
matrixC19_16,
matrixC19_17,
matrixC19_18,
matrixC19_19,
matrixC19_20,
matrixC19_21,
matrixC19_22,
matrixC19_23,
matrixC19_24,
matrixC19_25,
matrixC19_26,
matrixC19_27,
matrixC19_28,
matrixC19_29,
matrixC19_30,
matrixC19_31,
matrixC20_0,
matrixC20_1,
matrixC20_2,
matrixC20_3,
matrixC20_4,
matrixC20_5,
matrixC20_6,
matrixC20_7,
matrixC20_8,
matrixC20_9,
matrixC20_10,
matrixC20_11,
matrixC20_12,
matrixC20_13,
matrixC20_14,
matrixC20_15,
matrixC20_16,
matrixC20_17,
matrixC20_18,
matrixC20_19,
matrixC20_20,
matrixC20_21,
matrixC20_22,
matrixC20_23,
matrixC20_24,
matrixC20_25,
matrixC20_26,
matrixC20_27,
matrixC20_28,
matrixC20_29,
matrixC20_30,
matrixC20_31,
matrixC21_0,
matrixC21_1,
matrixC21_2,
matrixC21_3,
matrixC21_4,
matrixC21_5,
matrixC21_6,
matrixC21_7,
matrixC21_8,
matrixC21_9,
matrixC21_10,
matrixC21_11,
matrixC21_12,
matrixC21_13,
matrixC21_14,
matrixC21_15,
matrixC21_16,
matrixC21_17,
matrixC21_18,
matrixC21_19,
matrixC21_20,
matrixC21_21,
matrixC21_22,
matrixC21_23,
matrixC21_24,
matrixC21_25,
matrixC21_26,
matrixC21_27,
matrixC21_28,
matrixC21_29,
matrixC21_30,
matrixC21_31,
matrixC22_0,
matrixC22_1,
matrixC22_2,
matrixC22_3,
matrixC22_4,
matrixC22_5,
matrixC22_6,
matrixC22_7,
matrixC22_8,
matrixC22_9,
matrixC22_10,
matrixC22_11,
matrixC22_12,
matrixC22_13,
matrixC22_14,
matrixC22_15,
matrixC22_16,
matrixC22_17,
matrixC22_18,
matrixC22_19,
matrixC22_20,
matrixC22_21,
matrixC22_22,
matrixC22_23,
matrixC22_24,
matrixC22_25,
matrixC22_26,
matrixC22_27,
matrixC22_28,
matrixC22_29,
matrixC22_30,
matrixC22_31,
matrixC23_0,
matrixC23_1,
matrixC23_2,
matrixC23_3,
matrixC23_4,
matrixC23_5,
matrixC23_6,
matrixC23_7,
matrixC23_8,
matrixC23_9,
matrixC23_10,
matrixC23_11,
matrixC23_12,
matrixC23_13,
matrixC23_14,
matrixC23_15,
matrixC23_16,
matrixC23_17,
matrixC23_18,
matrixC23_19,
matrixC23_20,
matrixC23_21,
matrixC23_22,
matrixC23_23,
matrixC23_24,
matrixC23_25,
matrixC23_26,
matrixC23_27,
matrixC23_28,
matrixC23_29,
matrixC23_30,
matrixC23_31,
matrixC24_0,
matrixC24_1,
matrixC24_2,
matrixC24_3,
matrixC24_4,
matrixC24_5,
matrixC24_6,
matrixC24_7,
matrixC24_8,
matrixC24_9,
matrixC24_10,
matrixC24_11,
matrixC24_12,
matrixC24_13,
matrixC24_14,
matrixC24_15,
matrixC24_16,
matrixC24_17,
matrixC24_18,
matrixC24_19,
matrixC24_20,
matrixC24_21,
matrixC24_22,
matrixC24_23,
matrixC24_24,
matrixC24_25,
matrixC24_26,
matrixC24_27,
matrixC24_28,
matrixC24_29,
matrixC24_30,
matrixC24_31,
matrixC25_0,
matrixC25_1,
matrixC25_2,
matrixC25_3,
matrixC25_4,
matrixC25_5,
matrixC25_6,
matrixC25_7,
matrixC25_8,
matrixC25_9,
matrixC25_10,
matrixC25_11,
matrixC25_12,
matrixC25_13,
matrixC25_14,
matrixC25_15,
matrixC25_16,
matrixC25_17,
matrixC25_18,
matrixC25_19,
matrixC25_20,
matrixC25_21,
matrixC25_22,
matrixC25_23,
matrixC25_24,
matrixC25_25,
matrixC25_26,
matrixC25_27,
matrixC25_28,
matrixC25_29,
matrixC25_30,
matrixC25_31,
matrixC26_0,
matrixC26_1,
matrixC26_2,
matrixC26_3,
matrixC26_4,
matrixC26_5,
matrixC26_6,
matrixC26_7,
matrixC26_8,
matrixC26_9,
matrixC26_10,
matrixC26_11,
matrixC26_12,
matrixC26_13,
matrixC26_14,
matrixC26_15,
matrixC26_16,
matrixC26_17,
matrixC26_18,
matrixC26_19,
matrixC26_20,
matrixC26_21,
matrixC26_22,
matrixC26_23,
matrixC26_24,
matrixC26_25,
matrixC26_26,
matrixC26_27,
matrixC26_28,
matrixC26_29,
matrixC26_30,
matrixC26_31,
matrixC27_0,
matrixC27_1,
matrixC27_2,
matrixC27_3,
matrixC27_4,
matrixC27_5,
matrixC27_6,
matrixC27_7,
matrixC27_8,
matrixC27_9,
matrixC27_10,
matrixC27_11,
matrixC27_12,
matrixC27_13,
matrixC27_14,
matrixC27_15,
matrixC27_16,
matrixC27_17,
matrixC27_18,
matrixC27_19,
matrixC27_20,
matrixC27_21,
matrixC27_22,
matrixC27_23,
matrixC27_24,
matrixC27_25,
matrixC27_26,
matrixC27_27,
matrixC27_28,
matrixC27_29,
matrixC27_30,
matrixC27_31,
matrixC28_0,
matrixC28_1,
matrixC28_2,
matrixC28_3,
matrixC28_4,
matrixC28_5,
matrixC28_6,
matrixC28_7,
matrixC28_8,
matrixC28_9,
matrixC28_10,
matrixC28_11,
matrixC28_12,
matrixC28_13,
matrixC28_14,
matrixC28_15,
matrixC28_16,
matrixC28_17,
matrixC28_18,
matrixC28_19,
matrixC28_20,
matrixC28_21,
matrixC28_22,
matrixC28_23,
matrixC28_24,
matrixC28_25,
matrixC28_26,
matrixC28_27,
matrixC28_28,
matrixC28_29,
matrixC28_30,
matrixC28_31,
matrixC29_0,
matrixC29_1,
matrixC29_2,
matrixC29_3,
matrixC29_4,
matrixC29_5,
matrixC29_6,
matrixC29_7,
matrixC29_8,
matrixC29_9,
matrixC29_10,
matrixC29_11,
matrixC29_12,
matrixC29_13,
matrixC29_14,
matrixC29_15,
matrixC29_16,
matrixC29_17,
matrixC29_18,
matrixC29_19,
matrixC29_20,
matrixC29_21,
matrixC29_22,
matrixC29_23,
matrixC29_24,
matrixC29_25,
matrixC29_26,
matrixC29_27,
matrixC29_28,
matrixC29_29,
matrixC29_30,
matrixC29_31,
matrixC30_0,
matrixC30_1,
matrixC30_2,
matrixC30_3,
matrixC30_4,
matrixC30_5,
matrixC30_6,
matrixC30_7,
matrixC30_8,
matrixC30_9,
matrixC30_10,
matrixC30_11,
matrixC30_12,
matrixC30_13,
matrixC30_14,
matrixC30_15,
matrixC30_16,
matrixC30_17,
matrixC30_18,
matrixC30_19,
matrixC30_20,
matrixC30_21,
matrixC30_22,
matrixC30_23,
matrixC30_24,
matrixC30_25,
matrixC30_26,
matrixC30_27,
matrixC30_28,
matrixC30_29,
matrixC30_30,
matrixC30_31,
matrixC31_0,
matrixC31_1,
matrixC31_2,
matrixC31_3,
matrixC31_4,
matrixC31_5,
matrixC31_6,
matrixC31_7,
matrixC31_8,
matrixC31_9,
matrixC31_10,
matrixC31_11,
matrixC31_12,
matrixC31_13,
matrixC31_14,
matrixC31_15,
matrixC31_16,
matrixC31_17,
matrixC31_18,
matrixC31_19,
matrixC31_20,
matrixC31_21,
matrixC31_22,
matrixC31_23,
matrixC31_24,
matrixC31_25,
matrixC31_26,
matrixC31_27,
matrixC31_28,
matrixC31_29,
matrixC31_30,
matrixC31_31,

clk,
reset
);

input clk;
input reset;
input start_mat_mul;
input done_mat_mul;
input [`AWIDTH-1:0] address_mat_c;
input [`ADDR_STRIDE_WIDTH-1:0] address_stride_c;
input [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_in;
output [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out;
output [`AWIDTH-1:0] c_addr;
output c_data_available;
input [7:0] clk_cnt;
output row_latch_en;

input [7:0] final_mat_mul_size;
  input [`DWIDTH-1:0] matrixC0_0;
input [`DWIDTH-1:0] matrixC0_1;
input [`DWIDTH-1:0] matrixC0_2;
input [`DWIDTH-1:0] matrixC0_3;
input [`DWIDTH-1:0] matrixC0_4;
input [`DWIDTH-1:0] matrixC0_5;
input [`DWIDTH-1:0] matrixC0_6;
input [`DWIDTH-1:0] matrixC0_7;
input [`DWIDTH-1:0] matrixC0_8;
input [`DWIDTH-1:0] matrixC0_9;
input [`DWIDTH-1:0] matrixC0_10;
input [`DWIDTH-1:0] matrixC0_11;
input [`DWIDTH-1:0] matrixC0_12;
input [`DWIDTH-1:0] matrixC0_13;
input [`DWIDTH-1:0] matrixC0_14;
input [`DWIDTH-1:0] matrixC0_15;
input [`DWIDTH-1:0] matrixC0_16;
input [`DWIDTH-1:0] matrixC0_17;
input [`DWIDTH-1:0] matrixC0_18;
input [`DWIDTH-1:0] matrixC0_19;
input [`DWIDTH-1:0] matrixC0_20;
input [`DWIDTH-1:0] matrixC0_21;
input [`DWIDTH-1:0] matrixC0_22;
input [`DWIDTH-1:0] matrixC0_23;
input [`DWIDTH-1:0] matrixC0_24;
input [`DWIDTH-1:0] matrixC0_25;
input [`DWIDTH-1:0] matrixC0_26;
input [`DWIDTH-1:0] matrixC0_27;
input [`DWIDTH-1:0] matrixC0_28;
input [`DWIDTH-1:0] matrixC0_29;
input [`DWIDTH-1:0] matrixC0_30;
input [`DWIDTH-1:0] matrixC0_31;
input [`DWIDTH-1:0] matrixC1_0;
input [`DWIDTH-1:0] matrixC1_1;
input [`DWIDTH-1:0] matrixC1_2;
input [`DWIDTH-1:0] matrixC1_3;
input [`DWIDTH-1:0] matrixC1_4;
input [`DWIDTH-1:0] matrixC1_5;
input [`DWIDTH-1:0] matrixC1_6;
input [`DWIDTH-1:0] matrixC1_7;
input [`DWIDTH-1:0] matrixC1_8;
input [`DWIDTH-1:0] matrixC1_9;
input [`DWIDTH-1:0] matrixC1_10;
input [`DWIDTH-1:0] matrixC1_11;
input [`DWIDTH-1:0] matrixC1_12;
input [`DWIDTH-1:0] matrixC1_13;
input [`DWIDTH-1:0] matrixC1_14;
input [`DWIDTH-1:0] matrixC1_15;
input [`DWIDTH-1:0] matrixC1_16;
input [`DWIDTH-1:0] matrixC1_17;
input [`DWIDTH-1:0] matrixC1_18;
input [`DWIDTH-1:0] matrixC1_19;
input [`DWIDTH-1:0] matrixC1_20;
input [`DWIDTH-1:0] matrixC1_21;
input [`DWIDTH-1:0] matrixC1_22;
input [`DWIDTH-1:0] matrixC1_23;
input [`DWIDTH-1:0] matrixC1_24;
input [`DWIDTH-1:0] matrixC1_25;
input [`DWIDTH-1:0] matrixC1_26;
input [`DWIDTH-1:0] matrixC1_27;
input [`DWIDTH-1:0] matrixC1_28;
input [`DWIDTH-1:0] matrixC1_29;
input [`DWIDTH-1:0] matrixC1_30;
input [`DWIDTH-1:0] matrixC1_31;
input [`DWIDTH-1:0] matrixC2_0;
input [`DWIDTH-1:0] matrixC2_1;
input [`DWIDTH-1:0] matrixC2_2;
input [`DWIDTH-1:0] matrixC2_3;
input [`DWIDTH-1:0] matrixC2_4;
input [`DWIDTH-1:0] matrixC2_5;
input [`DWIDTH-1:0] matrixC2_6;
input [`DWIDTH-1:0] matrixC2_7;
input [`DWIDTH-1:0] matrixC2_8;
input [`DWIDTH-1:0] matrixC2_9;
input [`DWIDTH-1:0] matrixC2_10;
input [`DWIDTH-1:0] matrixC2_11;
input [`DWIDTH-1:0] matrixC2_12;
input [`DWIDTH-1:0] matrixC2_13;
input [`DWIDTH-1:0] matrixC2_14;
input [`DWIDTH-1:0] matrixC2_15;
input [`DWIDTH-1:0] matrixC2_16;
input [`DWIDTH-1:0] matrixC2_17;
input [`DWIDTH-1:0] matrixC2_18;
input [`DWIDTH-1:0] matrixC2_19;
input [`DWIDTH-1:0] matrixC2_20;
input [`DWIDTH-1:0] matrixC2_21;
input [`DWIDTH-1:0] matrixC2_22;
input [`DWIDTH-1:0] matrixC2_23;
input [`DWIDTH-1:0] matrixC2_24;
input [`DWIDTH-1:0] matrixC2_25;
input [`DWIDTH-1:0] matrixC2_26;
input [`DWIDTH-1:0] matrixC2_27;
input [`DWIDTH-1:0] matrixC2_28;
input [`DWIDTH-1:0] matrixC2_29;
input [`DWIDTH-1:0] matrixC2_30;
input [`DWIDTH-1:0] matrixC2_31;
input [`DWIDTH-1:0] matrixC3_0;
input [`DWIDTH-1:0] matrixC3_1;
input [`DWIDTH-1:0] matrixC3_2;
input [`DWIDTH-1:0] matrixC3_3;
input [`DWIDTH-1:0] matrixC3_4;
input [`DWIDTH-1:0] matrixC3_5;
input [`DWIDTH-1:0] matrixC3_6;
input [`DWIDTH-1:0] matrixC3_7;
input [`DWIDTH-1:0] matrixC3_8;
input [`DWIDTH-1:0] matrixC3_9;
input [`DWIDTH-1:0] matrixC3_10;
input [`DWIDTH-1:0] matrixC3_11;
input [`DWIDTH-1:0] matrixC3_12;
input [`DWIDTH-1:0] matrixC3_13;
input [`DWIDTH-1:0] matrixC3_14;
input [`DWIDTH-1:0] matrixC3_15;
input [`DWIDTH-1:0] matrixC3_16;
input [`DWIDTH-1:0] matrixC3_17;
input [`DWIDTH-1:0] matrixC3_18;
input [`DWIDTH-1:0] matrixC3_19;
input [`DWIDTH-1:0] matrixC3_20;
input [`DWIDTH-1:0] matrixC3_21;
input [`DWIDTH-1:0] matrixC3_22;
input [`DWIDTH-1:0] matrixC3_23;
input [`DWIDTH-1:0] matrixC3_24;
input [`DWIDTH-1:0] matrixC3_25;
input [`DWIDTH-1:0] matrixC3_26;
input [`DWIDTH-1:0] matrixC3_27;
input [`DWIDTH-1:0] matrixC3_28;
input [`DWIDTH-1:0] matrixC3_29;
input [`DWIDTH-1:0] matrixC3_30;
input [`DWIDTH-1:0] matrixC3_31;
input [`DWIDTH-1:0] matrixC4_0;
input [`DWIDTH-1:0] matrixC4_1;
input [`DWIDTH-1:0] matrixC4_2;
input [`DWIDTH-1:0] matrixC4_3;
input [`DWIDTH-1:0] matrixC4_4;
input [`DWIDTH-1:0] matrixC4_5;
input [`DWIDTH-1:0] matrixC4_6;
input [`DWIDTH-1:0] matrixC4_7;
input [`DWIDTH-1:0] matrixC4_8;
input [`DWIDTH-1:0] matrixC4_9;
input [`DWIDTH-1:0] matrixC4_10;
input [`DWIDTH-1:0] matrixC4_11;
input [`DWIDTH-1:0] matrixC4_12;
input [`DWIDTH-1:0] matrixC4_13;
input [`DWIDTH-1:0] matrixC4_14;
input [`DWIDTH-1:0] matrixC4_15;
input [`DWIDTH-1:0] matrixC4_16;
input [`DWIDTH-1:0] matrixC4_17;
input [`DWIDTH-1:0] matrixC4_18;
input [`DWIDTH-1:0] matrixC4_19;
input [`DWIDTH-1:0] matrixC4_20;
input [`DWIDTH-1:0] matrixC4_21;
input [`DWIDTH-1:0] matrixC4_22;
input [`DWIDTH-1:0] matrixC4_23;
input [`DWIDTH-1:0] matrixC4_24;
input [`DWIDTH-1:0] matrixC4_25;
input [`DWIDTH-1:0] matrixC4_26;
input [`DWIDTH-1:0] matrixC4_27;
input [`DWIDTH-1:0] matrixC4_28;
input [`DWIDTH-1:0] matrixC4_29;
input [`DWIDTH-1:0] matrixC4_30;
input [`DWIDTH-1:0] matrixC4_31;
input [`DWIDTH-1:0] matrixC5_0;
input [`DWIDTH-1:0] matrixC5_1;
input [`DWIDTH-1:0] matrixC5_2;
input [`DWIDTH-1:0] matrixC5_3;
input [`DWIDTH-1:0] matrixC5_4;
input [`DWIDTH-1:0] matrixC5_5;
input [`DWIDTH-1:0] matrixC5_6;
input [`DWIDTH-1:0] matrixC5_7;
input [`DWIDTH-1:0] matrixC5_8;
input [`DWIDTH-1:0] matrixC5_9;
input [`DWIDTH-1:0] matrixC5_10;
input [`DWIDTH-1:0] matrixC5_11;
input [`DWIDTH-1:0] matrixC5_12;
input [`DWIDTH-1:0] matrixC5_13;
input [`DWIDTH-1:0] matrixC5_14;
input [`DWIDTH-1:0] matrixC5_15;
input [`DWIDTH-1:0] matrixC5_16;
input [`DWIDTH-1:0] matrixC5_17;
input [`DWIDTH-1:0] matrixC5_18;
input [`DWIDTH-1:0] matrixC5_19;
input [`DWIDTH-1:0] matrixC5_20;
input [`DWIDTH-1:0] matrixC5_21;
input [`DWIDTH-1:0] matrixC5_22;
input [`DWIDTH-1:0] matrixC5_23;
input [`DWIDTH-1:0] matrixC5_24;
input [`DWIDTH-1:0] matrixC5_25;
input [`DWIDTH-1:0] matrixC5_26;
input [`DWIDTH-1:0] matrixC5_27;
input [`DWIDTH-1:0] matrixC5_28;
input [`DWIDTH-1:0] matrixC5_29;
input [`DWIDTH-1:0] matrixC5_30;
input [`DWIDTH-1:0] matrixC5_31;
input [`DWIDTH-1:0] matrixC6_0;
input [`DWIDTH-1:0] matrixC6_1;
input [`DWIDTH-1:0] matrixC6_2;
input [`DWIDTH-1:0] matrixC6_3;
input [`DWIDTH-1:0] matrixC6_4;
input [`DWIDTH-1:0] matrixC6_5;
input [`DWIDTH-1:0] matrixC6_6;
input [`DWIDTH-1:0] matrixC6_7;
input [`DWIDTH-1:0] matrixC6_8;
input [`DWIDTH-1:0] matrixC6_9;
input [`DWIDTH-1:0] matrixC6_10;
input [`DWIDTH-1:0] matrixC6_11;
input [`DWIDTH-1:0] matrixC6_12;
input [`DWIDTH-1:0] matrixC6_13;
input [`DWIDTH-1:0] matrixC6_14;
input [`DWIDTH-1:0] matrixC6_15;
input [`DWIDTH-1:0] matrixC6_16;
input [`DWIDTH-1:0] matrixC6_17;
input [`DWIDTH-1:0] matrixC6_18;
input [`DWIDTH-1:0] matrixC6_19;
input [`DWIDTH-1:0] matrixC6_20;
input [`DWIDTH-1:0] matrixC6_21;
input [`DWIDTH-1:0] matrixC6_22;
input [`DWIDTH-1:0] matrixC6_23;
input [`DWIDTH-1:0] matrixC6_24;
input [`DWIDTH-1:0] matrixC6_25;
input [`DWIDTH-1:0] matrixC6_26;
input [`DWIDTH-1:0] matrixC6_27;
input [`DWIDTH-1:0] matrixC6_28;
input [`DWIDTH-1:0] matrixC6_29;
input [`DWIDTH-1:0] matrixC6_30;
input [`DWIDTH-1:0] matrixC6_31;
input [`DWIDTH-1:0] matrixC7_0;
input [`DWIDTH-1:0] matrixC7_1;
input [`DWIDTH-1:0] matrixC7_2;
input [`DWIDTH-1:0] matrixC7_3;
input [`DWIDTH-1:0] matrixC7_4;
input [`DWIDTH-1:0] matrixC7_5;
input [`DWIDTH-1:0] matrixC7_6;
input [`DWIDTH-1:0] matrixC7_7;
input [`DWIDTH-1:0] matrixC7_8;
input [`DWIDTH-1:0] matrixC7_9;
input [`DWIDTH-1:0] matrixC7_10;
input [`DWIDTH-1:0] matrixC7_11;
input [`DWIDTH-1:0] matrixC7_12;
input [`DWIDTH-1:0] matrixC7_13;
input [`DWIDTH-1:0] matrixC7_14;
input [`DWIDTH-1:0] matrixC7_15;
input [`DWIDTH-1:0] matrixC7_16;
input [`DWIDTH-1:0] matrixC7_17;
input [`DWIDTH-1:0] matrixC7_18;
input [`DWIDTH-1:0] matrixC7_19;
input [`DWIDTH-1:0] matrixC7_20;
input [`DWIDTH-1:0] matrixC7_21;
input [`DWIDTH-1:0] matrixC7_22;
input [`DWIDTH-1:0] matrixC7_23;
input [`DWIDTH-1:0] matrixC7_24;
input [`DWIDTH-1:0] matrixC7_25;
input [`DWIDTH-1:0] matrixC7_26;
input [`DWIDTH-1:0] matrixC7_27;
input [`DWIDTH-1:0] matrixC7_28;
input [`DWIDTH-1:0] matrixC7_29;
input [`DWIDTH-1:0] matrixC7_30;
input [`DWIDTH-1:0] matrixC7_31;
input [`DWIDTH-1:0] matrixC8_0;
input [`DWIDTH-1:0] matrixC8_1;
input [`DWIDTH-1:0] matrixC8_2;
input [`DWIDTH-1:0] matrixC8_3;
input [`DWIDTH-1:0] matrixC8_4;
input [`DWIDTH-1:0] matrixC8_5;
input [`DWIDTH-1:0] matrixC8_6;
input [`DWIDTH-1:0] matrixC8_7;
input [`DWIDTH-1:0] matrixC8_8;
input [`DWIDTH-1:0] matrixC8_9;
input [`DWIDTH-1:0] matrixC8_10;
input [`DWIDTH-1:0] matrixC8_11;
input [`DWIDTH-1:0] matrixC8_12;
input [`DWIDTH-1:0] matrixC8_13;
input [`DWIDTH-1:0] matrixC8_14;
input [`DWIDTH-1:0] matrixC8_15;
input [`DWIDTH-1:0] matrixC8_16;
input [`DWIDTH-1:0] matrixC8_17;
input [`DWIDTH-1:0] matrixC8_18;
input [`DWIDTH-1:0] matrixC8_19;
input [`DWIDTH-1:0] matrixC8_20;
input [`DWIDTH-1:0] matrixC8_21;
input [`DWIDTH-1:0] matrixC8_22;
input [`DWIDTH-1:0] matrixC8_23;
input [`DWIDTH-1:0] matrixC8_24;
input [`DWIDTH-1:0] matrixC8_25;
input [`DWIDTH-1:0] matrixC8_26;
input [`DWIDTH-1:0] matrixC8_27;
input [`DWIDTH-1:0] matrixC8_28;
input [`DWIDTH-1:0] matrixC8_29;
input [`DWIDTH-1:0] matrixC8_30;
input [`DWIDTH-1:0] matrixC8_31;
input [`DWIDTH-1:0] matrixC9_0;
input [`DWIDTH-1:0] matrixC9_1;
input [`DWIDTH-1:0] matrixC9_2;
input [`DWIDTH-1:0] matrixC9_3;
input [`DWIDTH-1:0] matrixC9_4;
input [`DWIDTH-1:0] matrixC9_5;
input [`DWIDTH-1:0] matrixC9_6;
input [`DWIDTH-1:0] matrixC9_7;
input [`DWIDTH-1:0] matrixC9_8;
input [`DWIDTH-1:0] matrixC9_9;
input [`DWIDTH-1:0] matrixC9_10;
input [`DWIDTH-1:0] matrixC9_11;
input [`DWIDTH-1:0] matrixC9_12;
input [`DWIDTH-1:0] matrixC9_13;
input [`DWIDTH-1:0] matrixC9_14;
input [`DWIDTH-1:0] matrixC9_15;
input [`DWIDTH-1:0] matrixC9_16;
input [`DWIDTH-1:0] matrixC9_17;
input [`DWIDTH-1:0] matrixC9_18;
input [`DWIDTH-1:0] matrixC9_19;
input [`DWIDTH-1:0] matrixC9_20;
input [`DWIDTH-1:0] matrixC9_21;
input [`DWIDTH-1:0] matrixC9_22;
input [`DWIDTH-1:0] matrixC9_23;
input [`DWIDTH-1:0] matrixC9_24;
input [`DWIDTH-1:0] matrixC9_25;
input [`DWIDTH-1:0] matrixC9_26;
input [`DWIDTH-1:0] matrixC9_27;
input [`DWIDTH-1:0] matrixC9_28;
input [`DWIDTH-1:0] matrixC9_29;
input [`DWIDTH-1:0] matrixC9_30;
input [`DWIDTH-1:0] matrixC9_31;
input [`DWIDTH-1:0] matrixC10_0;
input [`DWIDTH-1:0] matrixC10_1;
input [`DWIDTH-1:0] matrixC10_2;
input [`DWIDTH-1:0] matrixC10_3;
input [`DWIDTH-1:0] matrixC10_4;
input [`DWIDTH-1:0] matrixC10_5;
input [`DWIDTH-1:0] matrixC10_6;
input [`DWIDTH-1:0] matrixC10_7;
input [`DWIDTH-1:0] matrixC10_8;
input [`DWIDTH-1:0] matrixC10_9;
input [`DWIDTH-1:0] matrixC10_10;
input [`DWIDTH-1:0] matrixC10_11;
input [`DWIDTH-1:0] matrixC10_12;
input [`DWIDTH-1:0] matrixC10_13;
input [`DWIDTH-1:0] matrixC10_14;
input [`DWIDTH-1:0] matrixC10_15;
input [`DWIDTH-1:0] matrixC10_16;
input [`DWIDTH-1:0] matrixC10_17;
input [`DWIDTH-1:0] matrixC10_18;
input [`DWIDTH-1:0] matrixC10_19;
input [`DWIDTH-1:0] matrixC10_20;
input [`DWIDTH-1:0] matrixC10_21;
input [`DWIDTH-1:0] matrixC10_22;
input [`DWIDTH-1:0] matrixC10_23;
input [`DWIDTH-1:0] matrixC10_24;
input [`DWIDTH-1:0] matrixC10_25;
input [`DWIDTH-1:0] matrixC10_26;
input [`DWIDTH-1:0] matrixC10_27;
input [`DWIDTH-1:0] matrixC10_28;
input [`DWIDTH-1:0] matrixC10_29;
input [`DWIDTH-1:0] matrixC10_30;
input [`DWIDTH-1:0] matrixC10_31;
input [`DWIDTH-1:0] matrixC11_0;
input [`DWIDTH-1:0] matrixC11_1;
input [`DWIDTH-1:0] matrixC11_2;
input [`DWIDTH-1:0] matrixC11_3;
input [`DWIDTH-1:0] matrixC11_4;
input [`DWIDTH-1:0] matrixC11_5;
input [`DWIDTH-1:0] matrixC11_6;
input [`DWIDTH-1:0] matrixC11_7;
input [`DWIDTH-1:0] matrixC11_8;
input [`DWIDTH-1:0] matrixC11_9;
input [`DWIDTH-1:0] matrixC11_10;
input [`DWIDTH-1:0] matrixC11_11;
input [`DWIDTH-1:0] matrixC11_12;
input [`DWIDTH-1:0] matrixC11_13;
input [`DWIDTH-1:0] matrixC11_14;
input [`DWIDTH-1:0] matrixC11_15;
input [`DWIDTH-1:0] matrixC11_16;
input [`DWIDTH-1:0] matrixC11_17;
input [`DWIDTH-1:0] matrixC11_18;
input [`DWIDTH-1:0] matrixC11_19;
input [`DWIDTH-1:0] matrixC11_20;
input [`DWIDTH-1:0] matrixC11_21;
input [`DWIDTH-1:0] matrixC11_22;
input [`DWIDTH-1:0] matrixC11_23;
input [`DWIDTH-1:0] matrixC11_24;
input [`DWIDTH-1:0] matrixC11_25;
input [`DWIDTH-1:0] matrixC11_26;
input [`DWIDTH-1:0] matrixC11_27;
input [`DWIDTH-1:0] matrixC11_28;
input [`DWIDTH-1:0] matrixC11_29;
input [`DWIDTH-1:0] matrixC11_30;
input [`DWIDTH-1:0] matrixC11_31;
input [`DWIDTH-1:0] matrixC12_0;
input [`DWIDTH-1:0] matrixC12_1;
input [`DWIDTH-1:0] matrixC12_2;
input [`DWIDTH-1:0] matrixC12_3;
input [`DWIDTH-1:0] matrixC12_4;
input [`DWIDTH-1:0] matrixC12_5;
input [`DWIDTH-1:0] matrixC12_6;
input [`DWIDTH-1:0] matrixC12_7;
input [`DWIDTH-1:0] matrixC12_8;
input [`DWIDTH-1:0] matrixC12_9;
input [`DWIDTH-1:0] matrixC12_10;
input [`DWIDTH-1:0] matrixC12_11;
input [`DWIDTH-1:0] matrixC12_12;
input [`DWIDTH-1:0] matrixC12_13;
input [`DWIDTH-1:0] matrixC12_14;
input [`DWIDTH-1:0] matrixC12_15;
input [`DWIDTH-1:0] matrixC12_16;
input [`DWIDTH-1:0] matrixC12_17;
input [`DWIDTH-1:0] matrixC12_18;
input [`DWIDTH-1:0] matrixC12_19;
input [`DWIDTH-1:0] matrixC12_20;
input [`DWIDTH-1:0] matrixC12_21;
input [`DWIDTH-1:0] matrixC12_22;
input [`DWIDTH-1:0] matrixC12_23;
input [`DWIDTH-1:0] matrixC12_24;
input [`DWIDTH-1:0] matrixC12_25;
input [`DWIDTH-1:0] matrixC12_26;
input [`DWIDTH-1:0] matrixC12_27;
input [`DWIDTH-1:0] matrixC12_28;
input [`DWIDTH-1:0] matrixC12_29;
input [`DWIDTH-1:0] matrixC12_30;
input [`DWIDTH-1:0] matrixC12_31;
input [`DWIDTH-1:0] matrixC13_0;
input [`DWIDTH-1:0] matrixC13_1;
input [`DWIDTH-1:0] matrixC13_2;
input [`DWIDTH-1:0] matrixC13_3;
input [`DWIDTH-1:0] matrixC13_4;
input [`DWIDTH-1:0] matrixC13_5;
input [`DWIDTH-1:0] matrixC13_6;
input [`DWIDTH-1:0] matrixC13_7;
input [`DWIDTH-1:0] matrixC13_8;
input [`DWIDTH-1:0] matrixC13_9;
input [`DWIDTH-1:0] matrixC13_10;
input [`DWIDTH-1:0] matrixC13_11;
input [`DWIDTH-1:0] matrixC13_12;
input [`DWIDTH-1:0] matrixC13_13;
input [`DWIDTH-1:0] matrixC13_14;
input [`DWIDTH-1:0] matrixC13_15;
input [`DWIDTH-1:0] matrixC13_16;
input [`DWIDTH-1:0] matrixC13_17;
input [`DWIDTH-1:0] matrixC13_18;
input [`DWIDTH-1:0] matrixC13_19;
input [`DWIDTH-1:0] matrixC13_20;
input [`DWIDTH-1:0] matrixC13_21;
input [`DWIDTH-1:0] matrixC13_22;
input [`DWIDTH-1:0] matrixC13_23;
input [`DWIDTH-1:0] matrixC13_24;
input [`DWIDTH-1:0] matrixC13_25;
input [`DWIDTH-1:0] matrixC13_26;
input [`DWIDTH-1:0] matrixC13_27;
input [`DWIDTH-1:0] matrixC13_28;
input [`DWIDTH-1:0] matrixC13_29;
input [`DWIDTH-1:0] matrixC13_30;
input [`DWIDTH-1:0] matrixC13_31;
input [`DWIDTH-1:0] matrixC14_0;
input [`DWIDTH-1:0] matrixC14_1;
input [`DWIDTH-1:0] matrixC14_2;
input [`DWIDTH-1:0] matrixC14_3;
input [`DWIDTH-1:0] matrixC14_4;
input [`DWIDTH-1:0] matrixC14_5;
input [`DWIDTH-1:0] matrixC14_6;
input [`DWIDTH-1:0] matrixC14_7;
input [`DWIDTH-1:0] matrixC14_8;
input [`DWIDTH-1:0] matrixC14_9;
input [`DWIDTH-1:0] matrixC14_10;
input [`DWIDTH-1:0] matrixC14_11;
input [`DWIDTH-1:0] matrixC14_12;
input [`DWIDTH-1:0] matrixC14_13;
input [`DWIDTH-1:0] matrixC14_14;
input [`DWIDTH-1:0] matrixC14_15;
input [`DWIDTH-1:0] matrixC14_16;
input [`DWIDTH-1:0] matrixC14_17;
input [`DWIDTH-1:0] matrixC14_18;
input [`DWIDTH-1:0] matrixC14_19;
input [`DWIDTH-1:0] matrixC14_20;
input [`DWIDTH-1:0] matrixC14_21;
input [`DWIDTH-1:0] matrixC14_22;
input [`DWIDTH-1:0] matrixC14_23;
input [`DWIDTH-1:0] matrixC14_24;
input [`DWIDTH-1:0] matrixC14_25;
input [`DWIDTH-1:0] matrixC14_26;
input [`DWIDTH-1:0] matrixC14_27;
input [`DWIDTH-1:0] matrixC14_28;
input [`DWIDTH-1:0] matrixC14_29;
input [`DWIDTH-1:0] matrixC14_30;
input [`DWIDTH-1:0] matrixC14_31;
input [`DWIDTH-1:0] matrixC15_0;
input [`DWIDTH-1:0] matrixC15_1;
input [`DWIDTH-1:0] matrixC15_2;
input [`DWIDTH-1:0] matrixC15_3;
input [`DWIDTH-1:0] matrixC15_4;
input [`DWIDTH-1:0] matrixC15_5;
input [`DWIDTH-1:0] matrixC15_6;
input [`DWIDTH-1:0] matrixC15_7;
input [`DWIDTH-1:0] matrixC15_8;
input [`DWIDTH-1:0] matrixC15_9;
input [`DWIDTH-1:0] matrixC15_10;
input [`DWIDTH-1:0] matrixC15_11;
input [`DWIDTH-1:0] matrixC15_12;
input [`DWIDTH-1:0] matrixC15_13;
input [`DWIDTH-1:0] matrixC15_14;
input [`DWIDTH-1:0] matrixC15_15;
input [`DWIDTH-1:0] matrixC15_16;
input [`DWIDTH-1:0] matrixC15_17;
input [`DWIDTH-1:0] matrixC15_18;
input [`DWIDTH-1:0] matrixC15_19;
input [`DWIDTH-1:0] matrixC15_20;
input [`DWIDTH-1:0] matrixC15_21;
input [`DWIDTH-1:0] matrixC15_22;
input [`DWIDTH-1:0] matrixC15_23;
input [`DWIDTH-1:0] matrixC15_24;
input [`DWIDTH-1:0] matrixC15_25;
input [`DWIDTH-1:0] matrixC15_26;
input [`DWIDTH-1:0] matrixC15_27;
input [`DWIDTH-1:0] matrixC15_28;
input [`DWIDTH-1:0] matrixC15_29;
input [`DWIDTH-1:0] matrixC15_30;
input [`DWIDTH-1:0] matrixC15_31;
input [`DWIDTH-1:0] matrixC16_0;
input [`DWIDTH-1:0] matrixC16_1;
input [`DWIDTH-1:0] matrixC16_2;
input [`DWIDTH-1:0] matrixC16_3;
input [`DWIDTH-1:0] matrixC16_4;
input [`DWIDTH-1:0] matrixC16_5;
input [`DWIDTH-1:0] matrixC16_6;
input [`DWIDTH-1:0] matrixC16_7;
input [`DWIDTH-1:0] matrixC16_8;
input [`DWIDTH-1:0] matrixC16_9;
input [`DWIDTH-1:0] matrixC16_10;
input [`DWIDTH-1:0] matrixC16_11;
input [`DWIDTH-1:0] matrixC16_12;
input [`DWIDTH-1:0] matrixC16_13;
input [`DWIDTH-1:0] matrixC16_14;
input [`DWIDTH-1:0] matrixC16_15;
input [`DWIDTH-1:0] matrixC16_16;
input [`DWIDTH-1:0] matrixC16_17;
input [`DWIDTH-1:0] matrixC16_18;
input [`DWIDTH-1:0] matrixC16_19;
input [`DWIDTH-1:0] matrixC16_20;
input [`DWIDTH-1:0] matrixC16_21;
input [`DWIDTH-1:0] matrixC16_22;
input [`DWIDTH-1:0] matrixC16_23;
input [`DWIDTH-1:0] matrixC16_24;
input [`DWIDTH-1:0] matrixC16_25;
input [`DWIDTH-1:0] matrixC16_26;
input [`DWIDTH-1:0] matrixC16_27;
input [`DWIDTH-1:0] matrixC16_28;
input [`DWIDTH-1:0] matrixC16_29;
input [`DWIDTH-1:0] matrixC16_30;
input [`DWIDTH-1:0] matrixC16_31;
input [`DWIDTH-1:0] matrixC17_0;
input [`DWIDTH-1:0] matrixC17_1;
input [`DWIDTH-1:0] matrixC17_2;
input [`DWIDTH-1:0] matrixC17_3;
input [`DWIDTH-1:0] matrixC17_4;
input [`DWIDTH-1:0] matrixC17_5;
input [`DWIDTH-1:0] matrixC17_6;
input [`DWIDTH-1:0] matrixC17_7;
input [`DWIDTH-1:0] matrixC17_8;
input [`DWIDTH-1:0] matrixC17_9;
input [`DWIDTH-1:0] matrixC17_10;
input [`DWIDTH-1:0] matrixC17_11;
input [`DWIDTH-1:0] matrixC17_12;
input [`DWIDTH-1:0] matrixC17_13;
input [`DWIDTH-1:0] matrixC17_14;
input [`DWIDTH-1:0] matrixC17_15;
input [`DWIDTH-1:0] matrixC17_16;
input [`DWIDTH-1:0] matrixC17_17;
input [`DWIDTH-1:0] matrixC17_18;
input [`DWIDTH-1:0] matrixC17_19;
input [`DWIDTH-1:0] matrixC17_20;
input [`DWIDTH-1:0] matrixC17_21;
input [`DWIDTH-1:0] matrixC17_22;
input [`DWIDTH-1:0] matrixC17_23;
input [`DWIDTH-1:0] matrixC17_24;
input [`DWIDTH-1:0] matrixC17_25;
input [`DWIDTH-1:0] matrixC17_26;
input [`DWIDTH-1:0] matrixC17_27;
input [`DWIDTH-1:0] matrixC17_28;
input [`DWIDTH-1:0] matrixC17_29;
input [`DWIDTH-1:0] matrixC17_30;
input [`DWIDTH-1:0] matrixC17_31;
input [`DWIDTH-1:0] matrixC18_0;
input [`DWIDTH-1:0] matrixC18_1;
input [`DWIDTH-1:0] matrixC18_2;
input [`DWIDTH-1:0] matrixC18_3;
input [`DWIDTH-1:0] matrixC18_4;
input [`DWIDTH-1:0] matrixC18_5;
input [`DWIDTH-1:0] matrixC18_6;
input [`DWIDTH-1:0] matrixC18_7;
input [`DWIDTH-1:0] matrixC18_8;
input [`DWIDTH-1:0] matrixC18_9;
input [`DWIDTH-1:0] matrixC18_10;
input [`DWIDTH-1:0] matrixC18_11;
input [`DWIDTH-1:0] matrixC18_12;
input [`DWIDTH-1:0] matrixC18_13;
input [`DWIDTH-1:0] matrixC18_14;
input [`DWIDTH-1:0] matrixC18_15;
input [`DWIDTH-1:0] matrixC18_16;
input [`DWIDTH-1:0] matrixC18_17;
input [`DWIDTH-1:0] matrixC18_18;
input [`DWIDTH-1:0] matrixC18_19;
input [`DWIDTH-1:0] matrixC18_20;
input [`DWIDTH-1:0] matrixC18_21;
input [`DWIDTH-1:0] matrixC18_22;
input [`DWIDTH-1:0] matrixC18_23;
input [`DWIDTH-1:0] matrixC18_24;
input [`DWIDTH-1:0] matrixC18_25;
input [`DWIDTH-1:0] matrixC18_26;
input [`DWIDTH-1:0] matrixC18_27;
input [`DWIDTH-1:0] matrixC18_28;
input [`DWIDTH-1:0] matrixC18_29;
input [`DWIDTH-1:0] matrixC18_30;
input [`DWIDTH-1:0] matrixC18_31;
input [`DWIDTH-1:0] matrixC19_0;
input [`DWIDTH-1:0] matrixC19_1;
input [`DWIDTH-1:0] matrixC19_2;
input [`DWIDTH-1:0] matrixC19_3;
input [`DWIDTH-1:0] matrixC19_4;
input [`DWIDTH-1:0] matrixC19_5;
input [`DWIDTH-1:0] matrixC19_6;
input [`DWIDTH-1:0] matrixC19_7;
input [`DWIDTH-1:0] matrixC19_8;
input [`DWIDTH-1:0] matrixC19_9;
input [`DWIDTH-1:0] matrixC19_10;
input [`DWIDTH-1:0] matrixC19_11;
input [`DWIDTH-1:0] matrixC19_12;
input [`DWIDTH-1:0] matrixC19_13;
input [`DWIDTH-1:0] matrixC19_14;
input [`DWIDTH-1:0] matrixC19_15;
input [`DWIDTH-1:0] matrixC19_16;
input [`DWIDTH-1:0] matrixC19_17;
input [`DWIDTH-1:0] matrixC19_18;
input [`DWIDTH-1:0] matrixC19_19;
input [`DWIDTH-1:0] matrixC19_20;
input [`DWIDTH-1:0] matrixC19_21;
input [`DWIDTH-1:0] matrixC19_22;
input [`DWIDTH-1:0] matrixC19_23;
input [`DWIDTH-1:0] matrixC19_24;
input [`DWIDTH-1:0] matrixC19_25;
input [`DWIDTH-1:0] matrixC19_26;
input [`DWIDTH-1:0] matrixC19_27;
input [`DWIDTH-1:0] matrixC19_28;
input [`DWIDTH-1:0] matrixC19_29;
input [`DWIDTH-1:0] matrixC19_30;
input [`DWIDTH-1:0] matrixC19_31;
input [`DWIDTH-1:0] matrixC20_0;
input [`DWIDTH-1:0] matrixC20_1;
input [`DWIDTH-1:0] matrixC20_2;
input [`DWIDTH-1:0] matrixC20_3;
input [`DWIDTH-1:0] matrixC20_4;
input [`DWIDTH-1:0] matrixC20_5;
input [`DWIDTH-1:0] matrixC20_6;
input [`DWIDTH-1:0] matrixC20_7;
input [`DWIDTH-1:0] matrixC20_8;
input [`DWIDTH-1:0] matrixC20_9;
input [`DWIDTH-1:0] matrixC20_10;
input [`DWIDTH-1:0] matrixC20_11;
input [`DWIDTH-1:0] matrixC20_12;
input [`DWIDTH-1:0] matrixC20_13;
input [`DWIDTH-1:0] matrixC20_14;
input [`DWIDTH-1:0] matrixC20_15;
input [`DWIDTH-1:0] matrixC20_16;
input [`DWIDTH-1:0] matrixC20_17;
input [`DWIDTH-1:0] matrixC20_18;
input [`DWIDTH-1:0] matrixC20_19;
input [`DWIDTH-1:0] matrixC20_20;
input [`DWIDTH-1:0] matrixC20_21;
input [`DWIDTH-1:0] matrixC20_22;
input [`DWIDTH-1:0] matrixC20_23;
input [`DWIDTH-1:0] matrixC20_24;
input [`DWIDTH-1:0] matrixC20_25;
input [`DWIDTH-1:0] matrixC20_26;
input [`DWIDTH-1:0] matrixC20_27;
input [`DWIDTH-1:0] matrixC20_28;
input [`DWIDTH-1:0] matrixC20_29;
input [`DWIDTH-1:0] matrixC20_30;
input [`DWIDTH-1:0] matrixC20_31;
input [`DWIDTH-1:0] matrixC21_0;
input [`DWIDTH-1:0] matrixC21_1;
input [`DWIDTH-1:0] matrixC21_2;
input [`DWIDTH-1:0] matrixC21_3;
input [`DWIDTH-1:0] matrixC21_4;
input [`DWIDTH-1:0] matrixC21_5;
input [`DWIDTH-1:0] matrixC21_6;
input [`DWIDTH-1:0] matrixC21_7;
input [`DWIDTH-1:0] matrixC21_8;
input [`DWIDTH-1:0] matrixC21_9;
input [`DWIDTH-1:0] matrixC21_10;
input [`DWIDTH-1:0] matrixC21_11;
input [`DWIDTH-1:0] matrixC21_12;
input [`DWIDTH-1:0] matrixC21_13;
input [`DWIDTH-1:0] matrixC21_14;
input [`DWIDTH-1:0] matrixC21_15;
input [`DWIDTH-1:0] matrixC21_16;
input [`DWIDTH-1:0] matrixC21_17;
input [`DWIDTH-1:0] matrixC21_18;
input [`DWIDTH-1:0] matrixC21_19;
input [`DWIDTH-1:0] matrixC21_20;
input [`DWIDTH-1:0] matrixC21_21;
input [`DWIDTH-1:0] matrixC21_22;
input [`DWIDTH-1:0] matrixC21_23;
input [`DWIDTH-1:0] matrixC21_24;
input [`DWIDTH-1:0] matrixC21_25;
input [`DWIDTH-1:0] matrixC21_26;
input [`DWIDTH-1:0] matrixC21_27;
input [`DWIDTH-1:0] matrixC21_28;
input [`DWIDTH-1:0] matrixC21_29;
input [`DWIDTH-1:0] matrixC21_30;
input [`DWIDTH-1:0] matrixC21_31;
input [`DWIDTH-1:0] matrixC22_0;
input [`DWIDTH-1:0] matrixC22_1;
input [`DWIDTH-1:0] matrixC22_2;
input [`DWIDTH-1:0] matrixC22_3;
input [`DWIDTH-1:0] matrixC22_4;
input [`DWIDTH-1:0] matrixC22_5;
input [`DWIDTH-1:0] matrixC22_6;
input [`DWIDTH-1:0] matrixC22_7;
input [`DWIDTH-1:0] matrixC22_8;
input [`DWIDTH-1:0] matrixC22_9;
input [`DWIDTH-1:0] matrixC22_10;
input [`DWIDTH-1:0] matrixC22_11;
input [`DWIDTH-1:0] matrixC22_12;
input [`DWIDTH-1:0] matrixC22_13;
input [`DWIDTH-1:0] matrixC22_14;
input [`DWIDTH-1:0] matrixC22_15;
input [`DWIDTH-1:0] matrixC22_16;
input [`DWIDTH-1:0] matrixC22_17;
input [`DWIDTH-1:0] matrixC22_18;
input [`DWIDTH-1:0] matrixC22_19;
input [`DWIDTH-1:0] matrixC22_20;
input [`DWIDTH-1:0] matrixC22_21;
input [`DWIDTH-1:0] matrixC22_22;
input [`DWIDTH-1:0] matrixC22_23;
input [`DWIDTH-1:0] matrixC22_24;
input [`DWIDTH-1:0] matrixC22_25;
input [`DWIDTH-1:0] matrixC22_26;
input [`DWIDTH-1:0] matrixC22_27;
input [`DWIDTH-1:0] matrixC22_28;
input [`DWIDTH-1:0] matrixC22_29;
input [`DWIDTH-1:0] matrixC22_30;
input [`DWIDTH-1:0] matrixC22_31;
input [`DWIDTH-1:0] matrixC23_0;
input [`DWIDTH-1:0] matrixC23_1;
input [`DWIDTH-1:0] matrixC23_2;
input [`DWIDTH-1:0] matrixC23_3;
input [`DWIDTH-1:0] matrixC23_4;
input [`DWIDTH-1:0] matrixC23_5;
input [`DWIDTH-1:0] matrixC23_6;
input [`DWIDTH-1:0] matrixC23_7;
input [`DWIDTH-1:0] matrixC23_8;
input [`DWIDTH-1:0] matrixC23_9;
input [`DWIDTH-1:0] matrixC23_10;
input [`DWIDTH-1:0] matrixC23_11;
input [`DWIDTH-1:0] matrixC23_12;
input [`DWIDTH-1:0] matrixC23_13;
input [`DWIDTH-1:0] matrixC23_14;
input [`DWIDTH-1:0] matrixC23_15;
input [`DWIDTH-1:0] matrixC23_16;
input [`DWIDTH-1:0] matrixC23_17;
input [`DWIDTH-1:0] matrixC23_18;
input [`DWIDTH-1:0] matrixC23_19;
input [`DWIDTH-1:0] matrixC23_20;
input [`DWIDTH-1:0] matrixC23_21;
input [`DWIDTH-1:0] matrixC23_22;
input [`DWIDTH-1:0] matrixC23_23;
input [`DWIDTH-1:0] matrixC23_24;
input [`DWIDTH-1:0] matrixC23_25;
input [`DWIDTH-1:0] matrixC23_26;
input [`DWIDTH-1:0] matrixC23_27;
input [`DWIDTH-1:0] matrixC23_28;
input [`DWIDTH-1:0] matrixC23_29;
input [`DWIDTH-1:0] matrixC23_30;
input [`DWIDTH-1:0] matrixC23_31;
input [`DWIDTH-1:0] matrixC24_0;
input [`DWIDTH-1:0] matrixC24_1;
input [`DWIDTH-1:0] matrixC24_2;
input [`DWIDTH-1:0] matrixC24_3;
input [`DWIDTH-1:0] matrixC24_4;
input [`DWIDTH-1:0] matrixC24_5;
input [`DWIDTH-1:0] matrixC24_6;
input [`DWIDTH-1:0] matrixC24_7;
input [`DWIDTH-1:0] matrixC24_8;
input [`DWIDTH-1:0] matrixC24_9;
input [`DWIDTH-1:0] matrixC24_10;
input [`DWIDTH-1:0] matrixC24_11;
input [`DWIDTH-1:0] matrixC24_12;
input [`DWIDTH-1:0] matrixC24_13;
input [`DWIDTH-1:0] matrixC24_14;
input [`DWIDTH-1:0] matrixC24_15;
input [`DWIDTH-1:0] matrixC24_16;
input [`DWIDTH-1:0] matrixC24_17;
input [`DWIDTH-1:0] matrixC24_18;
input [`DWIDTH-1:0] matrixC24_19;
input [`DWIDTH-1:0] matrixC24_20;
input [`DWIDTH-1:0] matrixC24_21;
input [`DWIDTH-1:0] matrixC24_22;
input [`DWIDTH-1:0] matrixC24_23;
input [`DWIDTH-1:0] matrixC24_24;
input [`DWIDTH-1:0] matrixC24_25;
input [`DWIDTH-1:0] matrixC24_26;
input [`DWIDTH-1:0] matrixC24_27;
input [`DWIDTH-1:0] matrixC24_28;
input [`DWIDTH-1:0] matrixC24_29;
input [`DWIDTH-1:0] matrixC24_30;
input [`DWIDTH-1:0] matrixC24_31;
input [`DWIDTH-1:0] matrixC25_0;
input [`DWIDTH-1:0] matrixC25_1;
input [`DWIDTH-1:0] matrixC25_2;
input [`DWIDTH-1:0] matrixC25_3;
input [`DWIDTH-1:0] matrixC25_4;
input [`DWIDTH-1:0] matrixC25_5;
input [`DWIDTH-1:0] matrixC25_6;
input [`DWIDTH-1:0] matrixC25_7;
input [`DWIDTH-1:0] matrixC25_8;
input [`DWIDTH-1:0] matrixC25_9;
input [`DWIDTH-1:0] matrixC25_10;
input [`DWIDTH-1:0] matrixC25_11;
input [`DWIDTH-1:0] matrixC25_12;
input [`DWIDTH-1:0] matrixC25_13;
input [`DWIDTH-1:0] matrixC25_14;
input [`DWIDTH-1:0] matrixC25_15;
input [`DWIDTH-1:0] matrixC25_16;
input [`DWIDTH-1:0] matrixC25_17;
input [`DWIDTH-1:0] matrixC25_18;
input [`DWIDTH-1:0] matrixC25_19;
input [`DWIDTH-1:0] matrixC25_20;
input [`DWIDTH-1:0] matrixC25_21;
input [`DWIDTH-1:0] matrixC25_22;
input [`DWIDTH-1:0] matrixC25_23;
input [`DWIDTH-1:0] matrixC25_24;
input [`DWIDTH-1:0] matrixC25_25;
input [`DWIDTH-1:0] matrixC25_26;
input [`DWIDTH-1:0] matrixC25_27;
input [`DWIDTH-1:0] matrixC25_28;
input [`DWIDTH-1:0] matrixC25_29;
input [`DWIDTH-1:0] matrixC25_30;
input [`DWIDTH-1:0] matrixC25_31;
input [`DWIDTH-1:0] matrixC26_0;
input [`DWIDTH-1:0] matrixC26_1;
input [`DWIDTH-1:0] matrixC26_2;
input [`DWIDTH-1:0] matrixC26_3;
input [`DWIDTH-1:0] matrixC26_4;
input [`DWIDTH-1:0] matrixC26_5;
input [`DWIDTH-1:0] matrixC26_6;
input [`DWIDTH-1:0] matrixC26_7;
input [`DWIDTH-1:0] matrixC26_8;
input [`DWIDTH-1:0] matrixC26_9;
input [`DWIDTH-1:0] matrixC26_10;
input [`DWIDTH-1:0] matrixC26_11;
input [`DWIDTH-1:0] matrixC26_12;
input [`DWIDTH-1:0] matrixC26_13;
input [`DWIDTH-1:0] matrixC26_14;
input [`DWIDTH-1:0] matrixC26_15;
input [`DWIDTH-1:0] matrixC26_16;
input [`DWIDTH-1:0] matrixC26_17;
input [`DWIDTH-1:0] matrixC26_18;
input [`DWIDTH-1:0] matrixC26_19;
input [`DWIDTH-1:0] matrixC26_20;
input [`DWIDTH-1:0] matrixC26_21;
input [`DWIDTH-1:0] matrixC26_22;
input [`DWIDTH-1:0] matrixC26_23;
input [`DWIDTH-1:0] matrixC26_24;
input [`DWIDTH-1:0] matrixC26_25;
input [`DWIDTH-1:0] matrixC26_26;
input [`DWIDTH-1:0] matrixC26_27;
input [`DWIDTH-1:0] matrixC26_28;
input [`DWIDTH-1:0] matrixC26_29;
input [`DWIDTH-1:0] matrixC26_30;
input [`DWIDTH-1:0] matrixC26_31;
input [`DWIDTH-1:0] matrixC27_0;
input [`DWIDTH-1:0] matrixC27_1;
input [`DWIDTH-1:0] matrixC27_2;
input [`DWIDTH-1:0] matrixC27_3;
input [`DWIDTH-1:0] matrixC27_4;
input [`DWIDTH-1:0] matrixC27_5;
input [`DWIDTH-1:0] matrixC27_6;
input [`DWIDTH-1:0] matrixC27_7;
input [`DWIDTH-1:0] matrixC27_8;
input [`DWIDTH-1:0] matrixC27_9;
input [`DWIDTH-1:0] matrixC27_10;
input [`DWIDTH-1:0] matrixC27_11;
input [`DWIDTH-1:0] matrixC27_12;
input [`DWIDTH-1:0] matrixC27_13;
input [`DWIDTH-1:0] matrixC27_14;
input [`DWIDTH-1:0] matrixC27_15;
input [`DWIDTH-1:0] matrixC27_16;
input [`DWIDTH-1:0] matrixC27_17;
input [`DWIDTH-1:0] matrixC27_18;
input [`DWIDTH-1:0] matrixC27_19;
input [`DWIDTH-1:0] matrixC27_20;
input [`DWIDTH-1:0] matrixC27_21;
input [`DWIDTH-1:0] matrixC27_22;
input [`DWIDTH-1:0] matrixC27_23;
input [`DWIDTH-1:0] matrixC27_24;
input [`DWIDTH-1:0] matrixC27_25;
input [`DWIDTH-1:0] matrixC27_26;
input [`DWIDTH-1:0] matrixC27_27;
input [`DWIDTH-1:0] matrixC27_28;
input [`DWIDTH-1:0] matrixC27_29;
input [`DWIDTH-1:0] matrixC27_30;
input [`DWIDTH-1:0] matrixC27_31;
input [`DWIDTH-1:0] matrixC28_0;
input [`DWIDTH-1:0] matrixC28_1;
input [`DWIDTH-1:0] matrixC28_2;
input [`DWIDTH-1:0] matrixC28_3;
input [`DWIDTH-1:0] matrixC28_4;
input [`DWIDTH-1:0] matrixC28_5;
input [`DWIDTH-1:0] matrixC28_6;
input [`DWIDTH-1:0] matrixC28_7;
input [`DWIDTH-1:0] matrixC28_8;
input [`DWIDTH-1:0] matrixC28_9;
input [`DWIDTH-1:0] matrixC28_10;
input [`DWIDTH-1:0] matrixC28_11;
input [`DWIDTH-1:0] matrixC28_12;
input [`DWIDTH-1:0] matrixC28_13;
input [`DWIDTH-1:0] matrixC28_14;
input [`DWIDTH-1:0] matrixC28_15;
input [`DWIDTH-1:0] matrixC28_16;
input [`DWIDTH-1:0] matrixC28_17;
input [`DWIDTH-1:0] matrixC28_18;
input [`DWIDTH-1:0] matrixC28_19;
input [`DWIDTH-1:0] matrixC28_20;
input [`DWIDTH-1:0] matrixC28_21;
input [`DWIDTH-1:0] matrixC28_22;
input [`DWIDTH-1:0] matrixC28_23;
input [`DWIDTH-1:0] matrixC28_24;
input [`DWIDTH-1:0] matrixC28_25;
input [`DWIDTH-1:0] matrixC28_26;
input [`DWIDTH-1:0] matrixC28_27;
input [`DWIDTH-1:0] matrixC28_28;
input [`DWIDTH-1:0] matrixC28_29;
input [`DWIDTH-1:0] matrixC28_30;
input [`DWIDTH-1:0] matrixC28_31;
input [`DWIDTH-1:0] matrixC29_0;
input [`DWIDTH-1:0] matrixC29_1;
input [`DWIDTH-1:0] matrixC29_2;
input [`DWIDTH-1:0] matrixC29_3;
input [`DWIDTH-1:0] matrixC29_4;
input [`DWIDTH-1:0] matrixC29_5;
input [`DWIDTH-1:0] matrixC29_6;
input [`DWIDTH-1:0] matrixC29_7;
input [`DWIDTH-1:0] matrixC29_8;
input [`DWIDTH-1:0] matrixC29_9;
input [`DWIDTH-1:0] matrixC29_10;
input [`DWIDTH-1:0] matrixC29_11;
input [`DWIDTH-1:0] matrixC29_12;
input [`DWIDTH-1:0] matrixC29_13;
input [`DWIDTH-1:0] matrixC29_14;
input [`DWIDTH-1:0] matrixC29_15;
input [`DWIDTH-1:0] matrixC29_16;
input [`DWIDTH-1:0] matrixC29_17;
input [`DWIDTH-1:0] matrixC29_18;
input [`DWIDTH-1:0] matrixC29_19;
input [`DWIDTH-1:0] matrixC29_20;
input [`DWIDTH-1:0] matrixC29_21;
input [`DWIDTH-1:0] matrixC29_22;
input [`DWIDTH-1:0] matrixC29_23;
input [`DWIDTH-1:0] matrixC29_24;
input [`DWIDTH-1:0] matrixC29_25;
input [`DWIDTH-1:0] matrixC29_26;
input [`DWIDTH-1:0] matrixC29_27;
input [`DWIDTH-1:0] matrixC29_28;
input [`DWIDTH-1:0] matrixC29_29;
input [`DWIDTH-1:0] matrixC29_30;
input [`DWIDTH-1:0] matrixC29_31;
input [`DWIDTH-1:0] matrixC30_0;
input [`DWIDTH-1:0] matrixC30_1;
input [`DWIDTH-1:0] matrixC30_2;
input [`DWIDTH-1:0] matrixC30_3;
input [`DWIDTH-1:0] matrixC30_4;
input [`DWIDTH-1:0] matrixC30_5;
input [`DWIDTH-1:0] matrixC30_6;
input [`DWIDTH-1:0] matrixC30_7;
input [`DWIDTH-1:0] matrixC30_8;
input [`DWIDTH-1:0] matrixC30_9;
input [`DWIDTH-1:0] matrixC30_10;
input [`DWIDTH-1:0] matrixC30_11;
input [`DWIDTH-1:0] matrixC30_12;
input [`DWIDTH-1:0] matrixC30_13;
input [`DWIDTH-1:0] matrixC30_14;
input [`DWIDTH-1:0] matrixC30_15;
input [`DWIDTH-1:0] matrixC30_16;
input [`DWIDTH-1:0] matrixC30_17;
input [`DWIDTH-1:0] matrixC30_18;
input [`DWIDTH-1:0] matrixC30_19;
input [`DWIDTH-1:0] matrixC30_20;
input [`DWIDTH-1:0] matrixC30_21;
input [`DWIDTH-1:0] matrixC30_22;
input [`DWIDTH-1:0] matrixC30_23;
input [`DWIDTH-1:0] matrixC30_24;
input [`DWIDTH-1:0] matrixC30_25;
input [`DWIDTH-1:0] matrixC30_26;
input [`DWIDTH-1:0] matrixC30_27;
input [`DWIDTH-1:0] matrixC30_28;
input [`DWIDTH-1:0] matrixC30_29;
input [`DWIDTH-1:0] matrixC30_30;
input [`DWIDTH-1:0] matrixC30_31;
input [`DWIDTH-1:0] matrixC31_0;
input [`DWIDTH-1:0] matrixC31_1;
input [`DWIDTH-1:0] matrixC31_2;
input [`DWIDTH-1:0] matrixC31_3;
input [`DWIDTH-1:0] matrixC31_4;
input [`DWIDTH-1:0] matrixC31_5;
input [`DWIDTH-1:0] matrixC31_6;
input [`DWIDTH-1:0] matrixC31_7;
input [`DWIDTH-1:0] matrixC31_8;
input [`DWIDTH-1:0] matrixC31_9;
input [`DWIDTH-1:0] matrixC31_10;
input [`DWIDTH-1:0] matrixC31_11;
input [`DWIDTH-1:0] matrixC31_12;
input [`DWIDTH-1:0] matrixC31_13;
input [`DWIDTH-1:0] matrixC31_14;
input [`DWIDTH-1:0] matrixC31_15;
input [`DWIDTH-1:0] matrixC31_16;
input [`DWIDTH-1:0] matrixC31_17;
input [`DWIDTH-1:0] matrixC31_18;
input [`DWIDTH-1:0] matrixC31_19;
input [`DWIDTH-1:0] matrixC31_20;
input [`DWIDTH-1:0] matrixC31_21;
input [`DWIDTH-1:0] matrixC31_22;
input [`DWIDTH-1:0] matrixC31_23;
input [`DWIDTH-1:0] matrixC31_24;
input [`DWIDTH-1:0] matrixC31_25;
input [`DWIDTH-1:0] matrixC31_26;
input [`DWIDTH-1:0] matrixC31_27;
input [`DWIDTH-1:0] matrixC31_28;
input [`DWIDTH-1:0] matrixC31_29;
input [`DWIDTH-1:0] matrixC31_30;
input [`DWIDTH-1:0] matrixC31_31;
wire row_latch_en;


//////////////////////////////////////////////////////////////////////////
// Logic to capture matrix C data from the PEs and shift it out
//////////////////////////////////////////////////////////////////////////
//assign row_latch_en = (clk_cnt==(`MAT_MUL_SIZE + (a_loc+b_loc) * `BB_MAT_MUL_SIZE + 10 +  `NUM_CYCLES_IN_MAC - 1));
//Writing the line above to avoid multiplication:
//assign row_latch_en = (clk_cnt==(`MAT_MUL_SIZE + ((a_loc+b_loc) << `LOG2_MAT_MUL_SIZE) + 10 +  `NUM_CYCLES_IN_MAC - 1));

assign row_latch_en =  
                       ((clk_cnt == ((final_mat_mul_size<<2) - final_mat_mul_size - 1 +`NUM_CYCLES_IN_MAC)));
    
reg c_data_available;
reg [`AWIDTH-1:0] c_addr;
reg start_capturing_c_data;
integer counter;
reg [32*`DWIDTH-1:0] c_data_out;
reg [32*`DWIDTH-1:0] c_data_out_1;
reg [32*`DWIDTH-1:0] c_data_out_2;
reg [32*`DWIDTH-1:0] c_data_out_3;
reg [32*`DWIDTH-1:0] c_data_out_4;
reg [32*`DWIDTH-1:0] c_data_out_5;
reg [32*`DWIDTH-1:0] c_data_out_6;
reg [32*`DWIDTH-1:0] c_data_out_7;
reg [32*`DWIDTH-1:0] c_data_out_8;
reg [32*`DWIDTH-1:0] c_data_out_9;
reg [32*`DWIDTH-1:0] c_data_out_10;
reg [32*`DWIDTH-1:0] c_data_out_11;
reg [32*`DWIDTH-1:0] c_data_out_12;
reg [32*`DWIDTH-1:0] c_data_out_13;
reg [32*`DWIDTH-1:0] c_data_out_14;
reg [32*`DWIDTH-1:0] c_data_out_15;
reg [32*`DWIDTH-1:0] c_data_out_16;
reg [32*`DWIDTH-1:0] c_data_out_17;
reg [32*`DWIDTH-1:0] c_data_out_18;
reg [32*`DWIDTH-1:0] c_data_out_19;
reg [32*`DWIDTH-1:0] c_data_out_20;
reg [32*`DWIDTH-1:0] c_data_out_21;
reg [32*`DWIDTH-1:0] c_data_out_22;
reg [32*`DWIDTH-1:0] c_data_out_23;
reg [32*`DWIDTH-1:0] c_data_out_24;
reg [32*`DWIDTH-1:0] c_data_out_25;
reg [32*`DWIDTH-1:0] c_data_out_26;
reg [32*`DWIDTH-1:0] c_data_out_27;
reg [32*`DWIDTH-1:0] c_data_out_28;
reg [32*`DWIDTH-1:0] c_data_out_29;
reg [32*`DWIDTH-1:0] c_data_out_30;
reg [32*`DWIDTH-1:0] c_data_out_31;
wire condition_to_start_shifting_output;
assign condition_to_start_shifting_output = 
                          row_latch_en ;  

  
//For larger matmuls, this logic will have more entries in the case statement
always @(posedge clk) begin
  if (reset | ~start_mat_mul) begin
    start_capturing_c_data <= 1'b0;
    c_data_available <= 1'b0;
    c_addr <= address_mat_c + address_stride_c;
    c_data_out <= 0;
    counter <= 0;

    c_data_out_1 <= 0;
    c_data_out_2 <= 0;
    c_data_out_3 <= 0;
    c_data_out_4 <= 0;
    c_data_out_5 <= 0;
    c_data_out_6 <= 0;
    c_data_out_7 <= 0;
    c_data_out_8 <= 0;
    c_data_out_9 <= 0;
    c_data_out_10 <= 0;
    c_data_out_11 <= 0;
    c_data_out_12 <= 0;
    c_data_out_13 <= 0;
    c_data_out_14 <= 0;
    c_data_out_15 <= 0;
    c_data_out_16 <= 0;
    c_data_out_17 <= 0;
    c_data_out_18 <= 0;
    c_data_out_19 <= 0;
    c_data_out_20 <= 0;
    c_data_out_21 <= 0;
    c_data_out_22 <= 0;
    c_data_out_23 <= 0;
    c_data_out_24 <= 0;
    c_data_out_25 <= 0;
    c_data_out_26 <= 0;
    c_data_out_27 <= 0;
    c_data_out_28 <= 0;
    c_data_out_29 <= 0;
    c_data_out_30 <= 0;
    c_data_out_31 <= 0;
  end else if (condition_to_start_shifting_output) begin
    start_capturing_c_data <= 1'b1;
    c_data_available <= 1'b1;
    c_addr <= c_addr - address_stride_c;
    c_data_out <= {matrixC31_31, matrixC30_31, matrixC29_31, matrixC28_31, matrixC27_31, matrixC26_31, matrixC25_31, matrixC24_31, matrixC23_31, matrixC22_31, matrixC21_31, matrixC20_31, matrixC19_31, matrixC18_31, matrixC17_31, matrixC16_31, matrixC15_31, matrixC14_31, matrixC13_31, matrixC12_31, matrixC11_31, matrixC10_31, matrixC9_31, matrixC8_31, matrixC7_31, matrixC6_31, matrixC5_31, matrixC4_31, matrixC3_31, matrixC2_31, matrixC1_31, matrixC0_31};
      c_data_out_1 <= {matrixC31_30, matrixC30_30, matrixC29_30, matrixC28_30, matrixC27_30, matrixC26_30, matrixC25_30, matrixC24_30, matrixC23_30, matrixC22_30, matrixC21_30, matrixC20_30, matrixC19_30, matrixC18_30, matrixC17_30, matrixC16_30, matrixC15_30, matrixC14_30, matrixC13_30, matrixC12_30, matrixC11_30, matrixC10_30, matrixC9_30, matrixC8_30, matrixC7_30, matrixC6_30, matrixC5_30, matrixC4_30, matrixC3_30, matrixC2_30, matrixC1_30, matrixC0_30};
      c_data_out_2 <= {matrixC31_29, matrixC30_29, matrixC29_29, matrixC28_29, matrixC27_29, matrixC26_29, matrixC25_29, matrixC24_29, matrixC23_29, matrixC22_29, matrixC21_29, matrixC20_29, matrixC19_29, matrixC18_29, matrixC17_29, matrixC16_29, matrixC15_29, matrixC14_29, matrixC13_29, matrixC12_29, matrixC11_29, matrixC10_29, matrixC9_29, matrixC8_29, matrixC7_29, matrixC6_29, matrixC5_29, matrixC4_29, matrixC3_29, matrixC2_29, matrixC1_29, matrixC0_29};
      c_data_out_3 <= {matrixC31_28, matrixC30_28, matrixC29_28, matrixC28_28, matrixC27_28, matrixC26_28, matrixC25_28, matrixC24_28, matrixC23_28, matrixC22_28, matrixC21_28, matrixC20_28, matrixC19_28, matrixC18_28, matrixC17_28, matrixC16_28, matrixC15_28, matrixC14_28, matrixC13_28, matrixC12_28, matrixC11_28, matrixC10_28, matrixC9_28, matrixC8_28, matrixC7_28, matrixC6_28, matrixC5_28, matrixC4_28, matrixC3_28, matrixC2_28, matrixC1_28, matrixC0_28};
      c_data_out_4 <= {matrixC31_27, matrixC30_27, matrixC29_27, matrixC28_27, matrixC27_27, matrixC26_27, matrixC25_27, matrixC24_27, matrixC23_27, matrixC22_27, matrixC21_27, matrixC20_27, matrixC19_27, matrixC18_27, matrixC17_27, matrixC16_27, matrixC15_27, matrixC14_27, matrixC13_27, matrixC12_27, matrixC11_27, matrixC10_27, matrixC9_27, matrixC8_27, matrixC7_27, matrixC6_27, matrixC5_27, matrixC4_27, matrixC3_27, matrixC2_27, matrixC1_27, matrixC0_27};
      c_data_out_5 <= {matrixC31_26, matrixC30_26, matrixC29_26, matrixC28_26, matrixC27_26, matrixC26_26, matrixC25_26, matrixC24_26, matrixC23_26, matrixC22_26, matrixC21_26, matrixC20_26, matrixC19_26, matrixC18_26, matrixC17_26, matrixC16_26, matrixC15_26, matrixC14_26, matrixC13_26, matrixC12_26, matrixC11_26, matrixC10_26, matrixC9_26, matrixC8_26, matrixC7_26, matrixC6_26, matrixC5_26, matrixC4_26, matrixC3_26, matrixC2_26, matrixC1_26, matrixC0_26};
      c_data_out_6 <= {matrixC31_25, matrixC30_25, matrixC29_25, matrixC28_25, matrixC27_25, matrixC26_25, matrixC25_25, matrixC24_25, matrixC23_25, matrixC22_25, matrixC21_25, matrixC20_25, matrixC19_25, matrixC18_25, matrixC17_25, matrixC16_25, matrixC15_25, matrixC14_25, matrixC13_25, matrixC12_25, matrixC11_25, matrixC10_25, matrixC9_25, matrixC8_25, matrixC7_25, matrixC6_25, matrixC5_25, matrixC4_25, matrixC3_25, matrixC2_25, matrixC1_25, matrixC0_25};
      c_data_out_7 <= {matrixC31_24, matrixC30_24, matrixC29_24, matrixC28_24, matrixC27_24, matrixC26_24, matrixC25_24, matrixC24_24, matrixC23_24, matrixC22_24, matrixC21_24, matrixC20_24, matrixC19_24, matrixC18_24, matrixC17_24, matrixC16_24, matrixC15_24, matrixC14_24, matrixC13_24, matrixC12_24, matrixC11_24, matrixC10_24, matrixC9_24, matrixC8_24, matrixC7_24, matrixC6_24, matrixC5_24, matrixC4_24, matrixC3_24, matrixC2_24, matrixC1_24, matrixC0_24};
      c_data_out_8 <= {matrixC31_23, matrixC30_23, matrixC29_23, matrixC28_23, matrixC27_23, matrixC26_23, matrixC25_23, matrixC24_23, matrixC23_23, matrixC22_23, matrixC21_23, matrixC20_23, matrixC19_23, matrixC18_23, matrixC17_23, matrixC16_23, matrixC15_23, matrixC14_23, matrixC13_23, matrixC12_23, matrixC11_23, matrixC10_23, matrixC9_23, matrixC8_23, matrixC7_23, matrixC6_23, matrixC5_23, matrixC4_23, matrixC3_23, matrixC2_23, matrixC1_23, matrixC0_23};
      c_data_out_9 <= {matrixC31_22, matrixC30_22, matrixC29_22, matrixC28_22, matrixC27_22, matrixC26_22, matrixC25_22, matrixC24_22, matrixC23_22, matrixC22_22, matrixC21_22, matrixC20_22, matrixC19_22, matrixC18_22, matrixC17_22, matrixC16_22, matrixC15_22, matrixC14_22, matrixC13_22, matrixC12_22, matrixC11_22, matrixC10_22, matrixC9_22, matrixC8_22, matrixC7_22, matrixC6_22, matrixC5_22, matrixC4_22, matrixC3_22, matrixC2_22, matrixC1_22, matrixC0_22};
      c_data_out_10 <= {matrixC31_21, matrixC30_21, matrixC29_21, matrixC28_21, matrixC27_21, matrixC26_21, matrixC25_21, matrixC24_21, matrixC23_21, matrixC22_21, matrixC21_21, matrixC20_21, matrixC19_21, matrixC18_21, matrixC17_21, matrixC16_21, matrixC15_21, matrixC14_21, matrixC13_21, matrixC12_21, matrixC11_21, matrixC10_21, matrixC9_21, matrixC8_21, matrixC7_21, matrixC6_21, matrixC5_21, matrixC4_21, matrixC3_21, matrixC2_21, matrixC1_21, matrixC0_21};
      c_data_out_11 <= {matrixC31_20, matrixC30_20, matrixC29_20, matrixC28_20, matrixC27_20, matrixC26_20, matrixC25_20, matrixC24_20, matrixC23_20, matrixC22_20, matrixC21_20, matrixC20_20, matrixC19_20, matrixC18_20, matrixC17_20, matrixC16_20, matrixC15_20, matrixC14_20, matrixC13_20, matrixC12_20, matrixC11_20, matrixC10_20, matrixC9_20, matrixC8_20, matrixC7_20, matrixC6_20, matrixC5_20, matrixC4_20, matrixC3_20, matrixC2_20, matrixC1_20, matrixC0_20};
      c_data_out_12 <= {matrixC31_19, matrixC30_19, matrixC29_19, matrixC28_19, matrixC27_19, matrixC26_19, matrixC25_19, matrixC24_19, matrixC23_19, matrixC22_19, matrixC21_19, matrixC20_19, matrixC19_19, matrixC18_19, matrixC17_19, matrixC16_19, matrixC15_19, matrixC14_19, matrixC13_19, matrixC12_19, matrixC11_19, matrixC10_19, matrixC9_19, matrixC8_19, matrixC7_19, matrixC6_19, matrixC5_19, matrixC4_19, matrixC3_19, matrixC2_19, matrixC1_19, matrixC0_19};
      c_data_out_13 <= {matrixC31_18, matrixC30_18, matrixC29_18, matrixC28_18, matrixC27_18, matrixC26_18, matrixC25_18, matrixC24_18, matrixC23_18, matrixC22_18, matrixC21_18, matrixC20_18, matrixC19_18, matrixC18_18, matrixC17_18, matrixC16_18, matrixC15_18, matrixC14_18, matrixC13_18, matrixC12_18, matrixC11_18, matrixC10_18, matrixC9_18, matrixC8_18, matrixC7_18, matrixC6_18, matrixC5_18, matrixC4_18, matrixC3_18, matrixC2_18, matrixC1_18, matrixC0_18};
      c_data_out_14 <= {matrixC31_17, matrixC30_17, matrixC29_17, matrixC28_17, matrixC27_17, matrixC26_17, matrixC25_17, matrixC24_17, matrixC23_17, matrixC22_17, matrixC21_17, matrixC20_17, matrixC19_17, matrixC18_17, matrixC17_17, matrixC16_17, matrixC15_17, matrixC14_17, matrixC13_17, matrixC12_17, matrixC11_17, matrixC10_17, matrixC9_17, matrixC8_17, matrixC7_17, matrixC6_17, matrixC5_17, matrixC4_17, matrixC3_17, matrixC2_17, matrixC1_17, matrixC0_17};
      c_data_out_15 <= {matrixC31_16, matrixC30_16, matrixC29_16, matrixC28_16, matrixC27_16, matrixC26_16, matrixC25_16, matrixC24_16, matrixC23_16, matrixC22_16, matrixC21_16, matrixC20_16, matrixC19_16, matrixC18_16, matrixC17_16, matrixC16_16, matrixC15_16, matrixC14_16, matrixC13_16, matrixC12_16, matrixC11_16, matrixC10_16, matrixC9_16, matrixC8_16, matrixC7_16, matrixC6_16, matrixC5_16, matrixC4_16, matrixC3_16, matrixC2_16, matrixC1_16, matrixC0_16};
      c_data_out_16 <= {matrixC31_15, matrixC30_15, matrixC29_15, matrixC28_15, matrixC27_15, matrixC26_15, matrixC25_15, matrixC24_15, matrixC23_15, matrixC22_15, matrixC21_15, matrixC20_15, matrixC19_15, matrixC18_15, matrixC17_15, matrixC16_15, matrixC15_15, matrixC14_15, matrixC13_15, matrixC12_15, matrixC11_15, matrixC10_15, matrixC9_15, matrixC8_15, matrixC7_15, matrixC6_15, matrixC5_15, matrixC4_15, matrixC3_15, matrixC2_15, matrixC1_15, matrixC0_15};
      c_data_out_17 <= {matrixC31_14, matrixC30_14, matrixC29_14, matrixC28_14, matrixC27_14, matrixC26_14, matrixC25_14, matrixC24_14, matrixC23_14, matrixC22_14, matrixC21_14, matrixC20_14, matrixC19_14, matrixC18_14, matrixC17_14, matrixC16_14, matrixC15_14, matrixC14_14, matrixC13_14, matrixC12_14, matrixC11_14, matrixC10_14, matrixC9_14, matrixC8_14, matrixC7_14, matrixC6_14, matrixC5_14, matrixC4_14, matrixC3_14, matrixC2_14, matrixC1_14, matrixC0_14};
      c_data_out_18 <= {matrixC31_13, matrixC30_13, matrixC29_13, matrixC28_13, matrixC27_13, matrixC26_13, matrixC25_13, matrixC24_13, matrixC23_13, matrixC22_13, matrixC21_13, matrixC20_13, matrixC19_13, matrixC18_13, matrixC17_13, matrixC16_13, matrixC15_13, matrixC14_13, matrixC13_13, matrixC12_13, matrixC11_13, matrixC10_13, matrixC9_13, matrixC8_13, matrixC7_13, matrixC6_13, matrixC5_13, matrixC4_13, matrixC3_13, matrixC2_13, matrixC1_13, matrixC0_13};
      c_data_out_19 <= {matrixC31_12, matrixC30_12, matrixC29_12, matrixC28_12, matrixC27_12, matrixC26_12, matrixC25_12, matrixC24_12, matrixC23_12, matrixC22_12, matrixC21_12, matrixC20_12, matrixC19_12, matrixC18_12, matrixC17_12, matrixC16_12, matrixC15_12, matrixC14_12, matrixC13_12, matrixC12_12, matrixC11_12, matrixC10_12, matrixC9_12, matrixC8_12, matrixC7_12, matrixC6_12, matrixC5_12, matrixC4_12, matrixC3_12, matrixC2_12, matrixC1_12, matrixC0_12};
      c_data_out_20 <= {matrixC31_11, matrixC30_11, matrixC29_11, matrixC28_11, matrixC27_11, matrixC26_11, matrixC25_11, matrixC24_11, matrixC23_11, matrixC22_11, matrixC21_11, matrixC20_11, matrixC19_11, matrixC18_11, matrixC17_11, matrixC16_11, matrixC15_11, matrixC14_11, matrixC13_11, matrixC12_11, matrixC11_11, matrixC10_11, matrixC9_11, matrixC8_11, matrixC7_11, matrixC6_11, matrixC5_11, matrixC4_11, matrixC3_11, matrixC2_11, matrixC1_11, matrixC0_11};
      c_data_out_21 <= {matrixC31_10, matrixC30_10, matrixC29_10, matrixC28_10, matrixC27_10, matrixC26_10, matrixC25_10, matrixC24_10, matrixC23_10, matrixC22_10, matrixC21_10, matrixC20_10, matrixC19_10, matrixC18_10, matrixC17_10, matrixC16_10, matrixC15_10, matrixC14_10, matrixC13_10, matrixC12_10, matrixC11_10, matrixC10_10, matrixC9_10, matrixC8_10, matrixC7_10, matrixC6_10, matrixC5_10, matrixC4_10, matrixC3_10, matrixC2_10, matrixC1_10, matrixC0_10};
      c_data_out_22 <= {matrixC31_9, matrixC30_9, matrixC29_9, matrixC28_9, matrixC27_9, matrixC26_9, matrixC25_9, matrixC24_9, matrixC23_9, matrixC22_9, matrixC21_9, matrixC20_9, matrixC19_9, matrixC18_9, matrixC17_9, matrixC16_9, matrixC15_9, matrixC14_9, matrixC13_9, matrixC12_9, matrixC11_9, matrixC10_9, matrixC9_9, matrixC8_9, matrixC7_9, matrixC6_9, matrixC5_9, matrixC4_9, matrixC3_9, matrixC2_9, matrixC1_9, matrixC0_9};
      c_data_out_23 <= {matrixC31_8, matrixC30_8, matrixC29_8, matrixC28_8, matrixC27_8, matrixC26_8, matrixC25_8, matrixC24_8, matrixC23_8, matrixC22_8, matrixC21_8, matrixC20_8, matrixC19_8, matrixC18_8, matrixC17_8, matrixC16_8, matrixC15_8, matrixC14_8, matrixC13_8, matrixC12_8, matrixC11_8, matrixC10_8, matrixC9_8, matrixC8_8, matrixC7_8, matrixC6_8, matrixC5_8, matrixC4_8, matrixC3_8, matrixC2_8, matrixC1_8, matrixC0_8};
      c_data_out_24 <= {matrixC31_7, matrixC30_7, matrixC29_7, matrixC28_7, matrixC27_7, matrixC26_7, matrixC25_7, matrixC24_7, matrixC23_7, matrixC22_7, matrixC21_7, matrixC20_7, matrixC19_7, matrixC18_7, matrixC17_7, matrixC16_7, matrixC15_7, matrixC14_7, matrixC13_7, matrixC12_7, matrixC11_7, matrixC10_7, matrixC9_7, matrixC8_7, matrixC7_7, matrixC6_7, matrixC5_7, matrixC4_7, matrixC3_7, matrixC2_7, matrixC1_7, matrixC0_7};
      c_data_out_25 <= {matrixC31_6, matrixC30_6, matrixC29_6, matrixC28_6, matrixC27_6, matrixC26_6, matrixC25_6, matrixC24_6, matrixC23_6, matrixC22_6, matrixC21_6, matrixC20_6, matrixC19_6, matrixC18_6, matrixC17_6, matrixC16_6, matrixC15_6, matrixC14_6, matrixC13_6, matrixC12_6, matrixC11_6, matrixC10_6, matrixC9_6, matrixC8_6, matrixC7_6, matrixC6_6, matrixC5_6, matrixC4_6, matrixC3_6, matrixC2_6, matrixC1_6, matrixC0_6};
      c_data_out_26 <= {matrixC31_5, matrixC30_5, matrixC29_5, matrixC28_5, matrixC27_5, matrixC26_5, matrixC25_5, matrixC24_5, matrixC23_5, matrixC22_5, matrixC21_5, matrixC20_5, matrixC19_5, matrixC18_5, matrixC17_5, matrixC16_5, matrixC15_5, matrixC14_5, matrixC13_5, matrixC12_5, matrixC11_5, matrixC10_5, matrixC9_5, matrixC8_5, matrixC7_5, matrixC6_5, matrixC5_5, matrixC4_5, matrixC3_5, matrixC2_5, matrixC1_5, matrixC0_5};
      c_data_out_27 <= {matrixC31_4, matrixC30_4, matrixC29_4, matrixC28_4, matrixC27_4, matrixC26_4, matrixC25_4, matrixC24_4, matrixC23_4, matrixC22_4, matrixC21_4, matrixC20_4, matrixC19_4, matrixC18_4, matrixC17_4, matrixC16_4, matrixC15_4, matrixC14_4, matrixC13_4, matrixC12_4, matrixC11_4, matrixC10_4, matrixC9_4, matrixC8_4, matrixC7_4, matrixC6_4, matrixC5_4, matrixC4_4, matrixC3_4, matrixC2_4, matrixC1_4, matrixC0_4};
      c_data_out_28 <= {matrixC31_3, matrixC30_3, matrixC29_3, matrixC28_3, matrixC27_3, matrixC26_3, matrixC25_3, matrixC24_3, matrixC23_3, matrixC22_3, matrixC21_3, matrixC20_3, matrixC19_3, matrixC18_3, matrixC17_3, matrixC16_3, matrixC15_3, matrixC14_3, matrixC13_3, matrixC12_3, matrixC11_3, matrixC10_3, matrixC9_3, matrixC8_3, matrixC7_3, matrixC6_3, matrixC5_3, matrixC4_3, matrixC3_3, matrixC2_3, matrixC1_3, matrixC0_3};
      c_data_out_29 <= {matrixC31_2, matrixC30_2, matrixC29_2, matrixC28_2, matrixC27_2, matrixC26_2, matrixC25_2, matrixC24_2, matrixC23_2, matrixC22_2, matrixC21_2, matrixC20_2, matrixC19_2, matrixC18_2, matrixC17_2, matrixC16_2, matrixC15_2, matrixC14_2, matrixC13_2, matrixC12_2, matrixC11_2, matrixC10_2, matrixC9_2, matrixC8_2, matrixC7_2, matrixC6_2, matrixC5_2, matrixC4_2, matrixC3_2, matrixC2_2, matrixC1_2, matrixC0_2};
      c_data_out_30 <= {matrixC31_1, matrixC30_1, matrixC29_1, matrixC28_1, matrixC27_1, matrixC26_1, matrixC25_1, matrixC24_1, matrixC23_1, matrixC22_1, matrixC21_1, matrixC20_1, matrixC19_1, matrixC18_1, matrixC17_1, matrixC16_1, matrixC15_1, matrixC14_1, matrixC13_1, matrixC12_1, matrixC11_1, matrixC10_1, matrixC9_1, matrixC8_1, matrixC7_1, matrixC6_1, matrixC5_1, matrixC4_1, matrixC3_1, matrixC2_1, matrixC1_1, matrixC0_1};
      c_data_out_31 <= {matrixC31_0, matrixC30_0, matrixC29_0, matrixC28_0, matrixC27_0, matrixC26_0, matrixC25_0, matrixC24_0, matrixC23_0, matrixC22_0, matrixC21_0, matrixC20_0, matrixC19_0, matrixC18_0, matrixC17_0, matrixC16_0, matrixC15_0, matrixC14_0, matrixC13_0, matrixC12_0, matrixC11_0, matrixC10_0, matrixC9_0, matrixC8_0, matrixC7_0, matrixC6_0, matrixC5_0, matrixC4_0, matrixC3_0, matrixC2_0, matrixC1_0, matrixC0_0};

    counter <= counter + 1;
  end else if (done_mat_mul) begin
    start_capturing_c_data <= 1'b0;
    c_data_available <= 1'b0;
    c_addr <= address_mat_c + address_stride_c;
    c_data_out <= 0;

    c_data_out_1 <= 0;
    c_data_out_2 <= 0;
    c_data_out_3 <= 0;
    c_data_out_4 <= 0;
    c_data_out_5 <= 0;
    c_data_out_6 <= 0;
    c_data_out_7 <= 0;
    c_data_out_8 <= 0;
    c_data_out_9 <= 0;
    c_data_out_10 <= 0;
    c_data_out_11 <= 0;
    c_data_out_12 <= 0;
    c_data_out_13 <= 0;
    c_data_out_14 <= 0;
    c_data_out_15 <= 0;
    c_data_out_16 <= 0;
    c_data_out_17 <= 0;
    c_data_out_18 <= 0;
    c_data_out_19 <= 0;
    c_data_out_20 <= 0;
    c_data_out_21 <= 0;
    c_data_out_22 <= 0;
    c_data_out_23 <= 0;
    c_data_out_24 <= 0;
    c_data_out_25 <= 0;
    c_data_out_26 <= 0;
    c_data_out_27 <= 0;
    c_data_out_28 <= 0;
    c_data_out_29 <= 0;
    c_data_out_30 <= 0;
    c_data_out_31 <= 0;
  end 
  else if (counter >= `MAT_MUL_SIZE) begin
    c_data_out <= c_data_out_1;
    c_addr <= c_addr - address_stride_c; 

    c_data_out_1 <= c_data_out_2;
    c_data_out_2 <= c_data_out_3;
    c_data_out_3 <= c_data_out_4;
    c_data_out_4 <= c_data_out_5;
    c_data_out_5 <= c_data_out_6;
    c_data_out_6 <= c_data_out_7;
    c_data_out_7 <= c_data_out_8;
    c_data_out_8 <= c_data_out_9;
    c_data_out_9 <= c_data_out_10;
    c_data_out_10 <= c_data_out_11;
    c_data_out_11 <= c_data_out_12;
    c_data_out_12 <= c_data_out_13;
    c_data_out_13 <= c_data_out_14;
    c_data_out_14 <= c_data_out_15;
    c_data_out_15 <= c_data_out_16;
    c_data_out_16 <= c_data_out_17;
    c_data_out_17 <= c_data_out_18;
    c_data_out_18 <= c_data_out_19;
    c_data_out_19 <= c_data_out_20;
    c_data_out_20 <= c_data_out_21;
    c_data_out_21 <= c_data_out_22;
    c_data_out_22 <= c_data_out_23;
    c_data_out_23 <= c_data_out_24;
    c_data_out_24 <= c_data_out_25;
    c_data_out_25 <= c_data_out_26;
    c_data_out_26 <= c_data_out_27;
    c_data_out_27 <= c_data_out_28;
    c_data_out_28 <= c_data_out_29;
    c_data_out_29 <= c_data_out_30;
    c_data_out_30 <= c_data_out_31;
    c_data_out_31 <= c_data_in;
  end
  else if (start_capturing_c_data) begin
    c_data_available <= 1'b1;
    c_addr <= c_addr - address_stride_c; 
    counter <= counter + 1;
    c_data_out <= c_data_out_1;

    c_data_out_1 <= c_data_out_2;
    c_data_out_2 <= c_data_out_3;
    c_data_out_3 <= c_data_out_4;
    c_data_out_4 <= c_data_out_5;
    c_data_out_5 <= c_data_out_6;
    c_data_out_6 <= c_data_out_7;
    c_data_out_7 <= c_data_out_8;
    c_data_out_8 <= c_data_out_9;
    c_data_out_9 <= c_data_out_10;
    c_data_out_10 <= c_data_out_11;
    c_data_out_11 <= c_data_out_12;
    c_data_out_12 <= c_data_out_13;
    c_data_out_13 <= c_data_out_14;
    c_data_out_14 <= c_data_out_15;
    c_data_out_15 <= c_data_out_16;
    c_data_out_16 <= c_data_out_17;
    c_data_out_17 <= c_data_out_18;
    c_data_out_18 <= c_data_out_19;
    c_data_out_19 <= c_data_out_20;
    c_data_out_20 <= c_data_out_21;
    c_data_out_21 <= c_data_out_22;
    c_data_out_22 <= c_data_out_23;
    c_data_out_23 <= c_data_out_24;
    c_data_out_24 <= c_data_out_25;
    c_data_out_25 <= c_data_out_26;
    c_data_out_26 <= c_data_out_27;
    c_data_out_27 <= c_data_out_28;
    c_data_out_28 <= c_data_out_29;
    c_data_out_29 <= c_data_out_30;
    c_data_out_30 <= c_data_out_31;
    c_data_out_31 <= c_data_in;
  end
end

endmodule


//////////////////////////////////////////////////////////////////////////
// Systolic data setup
//////////////////////////////////////////////////////////////////////////
module systolic_data_setup(
clk,
reset,
start_mat_mul,
a_addr,
b_addr,
address_mat_a,
address_mat_b,
address_stride_a,
address_stride_b,
a_data,
b_data,
clk_cnt,
a0_data,
b0_data,
a1_data_delayed_1,
b1_data_delayed_1,
a2_data_delayed_2,
b2_data_delayed_2,
a3_data_delayed_3,
b3_data_delayed_3,
a4_data_delayed_4,
b4_data_delayed_4,
a5_data_delayed_5,
b5_data_delayed_5,
a6_data_delayed_6,
b6_data_delayed_6,
a7_data_delayed_7,
b7_data_delayed_7,
a8_data_delayed_8,
b8_data_delayed_8,
a9_data_delayed_9,
b9_data_delayed_9,
a10_data_delayed_10,
b10_data_delayed_10,
a11_data_delayed_11,
b11_data_delayed_11,
a12_data_delayed_12,
b12_data_delayed_12,
a13_data_delayed_13,
b13_data_delayed_13,
a14_data_delayed_14,
b14_data_delayed_14,
a15_data_delayed_15,
b15_data_delayed_15,
a16_data_delayed_16,
b16_data_delayed_16,
a17_data_delayed_17,
b17_data_delayed_17,
a18_data_delayed_18,
b18_data_delayed_18,
a19_data_delayed_19,
b19_data_delayed_19,
a20_data_delayed_20,
b20_data_delayed_20,
a21_data_delayed_21,
b21_data_delayed_21,
a22_data_delayed_22,
b22_data_delayed_22,
a23_data_delayed_23,
b23_data_delayed_23,
a24_data_delayed_24,
b24_data_delayed_24,
a25_data_delayed_25,
b25_data_delayed_25,
a26_data_delayed_26,
b26_data_delayed_26,
a27_data_delayed_27,
b27_data_delayed_27,
a28_data_delayed_28,
b28_data_delayed_28,
a29_data_delayed_29,
b29_data_delayed_29,
a30_data_delayed_30,
b30_data_delayed_30,
a31_data_delayed_31,
b31_data_delayed_31,

validity_mask_a_rows,
validity_mask_a_cols_b_rows,
validity_mask_b_cols,

final_mat_mul_size,
  
a_loc,
b_loc
);

input clk;
input reset;
input start_mat_mul;
output [`AWIDTH-1:0] a_addr;
output [`AWIDTH-1:0] b_addr;
input [`AWIDTH-1:0] address_mat_a;
input [`AWIDTH-1:0] address_mat_b;
input [`ADDR_STRIDE_WIDTH-1:0] address_stride_a;
input [`ADDR_STRIDE_WIDTH-1:0] address_stride_b;
input [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data;
input [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data;
input [7:0] clk_cnt;
output [`DWIDTH-1:0] a0_data;
output [`DWIDTH-1:0] b0_data;
output [`DWIDTH-1:0] a1_data_delayed_1;
output [`DWIDTH-1:0] b1_data_delayed_1;
output [`DWIDTH-1:0] a2_data_delayed_2;
output [`DWIDTH-1:0] b2_data_delayed_2;
output [`DWIDTH-1:0] a3_data_delayed_3;
output [`DWIDTH-1:0] b3_data_delayed_3;
output [`DWIDTH-1:0] a4_data_delayed_4;
output [`DWIDTH-1:0] b4_data_delayed_4;
output [`DWIDTH-1:0] a5_data_delayed_5;
output [`DWIDTH-1:0] b5_data_delayed_5;
output [`DWIDTH-1:0] a6_data_delayed_6;
output [`DWIDTH-1:0] b6_data_delayed_6;
output [`DWIDTH-1:0] a7_data_delayed_7;
output [`DWIDTH-1:0] b7_data_delayed_7;
output [`DWIDTH-1:0] a8_data_delayed_8;
output [`DWIDTH-1:0] b8_data_delayed_8;
output [`DWIDTH-1:0] a9_data_delayed_9;
output [`DWIDTH-1:0] b9_data_delayed_9;
output [`DWIDTH-1:0] a10_data_delayed_10;
output [`DWIDTH-1:0] b10_data_delayed_10;
output [`DWIDTH-1:0] a11_data_delayed_11;
output [`DWIDTH-1:0] b11_data_delayed_11;
output [`DWIDTH-1:0] a12_data_delayed_12;
output [`DWIDTH-1:0] b12_data_delayed_12;
output [`DWIDTH-1:0] a13_data_delayed_13;
output [`DWIDTH-1:0] b13_data_delayed_13;
output [`DWIDTH-1:0] a14_data_delayed_14;
output [`DWIDTH-1:0] b14_data_delayed_14;
output [`DWIDTH-1:0] a15_data_delayed_15;
output [`DWIDTH-1:0] b15_data_delayed_15;
output [`DWIDTH-1:0] a16_data_delayed_16;
output [`DWIDTH-1:0] b16_data_delayed_16;
output [`DWIDTH-1:0] a17_data_delayed_17;
output [`DWIDTH-1:0] b17_data_delayed_17;
output [`DWIDTH-1:0] a18_data_delayed_18;
output [`DWIDTH-1:0] b18_data_delayed_18;
output [`DWIDTH-1:0] a19_data_delayed_19;
output [`DWIDTH-1:0] b19_data_delayed_19;
output [`DWIDTH-1:0] a20_data_delayed_20;
output [`DWIDTH-1:0] b20_data_delayed_20;
output [`DWIDTH-1:0] a21_data_delayed_21;
output [`DWIDTH-1:0] b21_data_delayed_21;
output [`DWIDTH-1:0] a22_data_delayed_22;
output [`DWIDTH-1:0] b22_data_delayed_22;
output [`DWIDTH-1:0] a23_data_delayed_23;
output [`DWIDTH-1:0] b23_data_delayed_23;
output [`DWIDTH-1:0] a24_data_delayed_24;
output [`DWIDTH-1:0] b24_data_delayed_24;
output [`DWIDTH-1:0] a25_data_delayed_25;
output [`DWIDTH-1:0] b25_data_delayed_25;
output [`DWIDTH-1:0] a26_data_delayed_26;
output [`DWIDTH-1:0] b26_data_delayed_26;
output [`DWIDTH-1:0] a27_data_delayed_27;
output [`DWIDTH-1:0] b27_data_delayed_27;
output [`DWIDTH-1:0] a28_data_delayed_28;
output [`DWIDTH-1:0] b28_data_delayed_28;
output [`DWIDTH-1:0] a29_data_delayed_29;
output [`DWIDTH-1:0] b29_data_delayed_29;
output [`DWIDTH-1:0] a30_data_delayed_30;
output [`DWIDTH-1:0] b30_data_delayed_30;
output [`DWIDTH-1:0] a31_data_delayed_31;
output [`DWIDTH-1:0] b31_data_delayed_31;

input [`MASK_WIDTH-1:0] validity_mask_a_rows;
input [`MASK_WIDTH-1:0] validity_mask_a_cols_b_rows;
input [`MASK_WIDTH-1:0] validity_mask_b_cols;

input [7:0] final_mat_mul_size;
  
input [7:0] a_loc;
input [7:0] b_loc;
wire [`DWIDTH-1:0] a0_data;
wire [`DWIDTH-1:0] a1_data;
wire [`DWIDTH-1:0] a2_data;
wire [`DWIDTH-1:0] a3_data;
wire [`DWIDTH-1:0] a4_data;
wire [`DWIDTH-1:0] a5_data;
wire [`DWIDTH-1:0] a6_data;
wire [`DWIDTH-1:0] a7_data;
wire [`DWIDTH-1:0] a8_data;
wire [`DWIDTH-1:0] a9_data;
wire [`DWIDTH-1:0] a10_data;
wire [`DWIDTH-1:0] a11_data;
wire [`DWIDTH-1:0] a12_data;
wire [`DWIDTH-1:0] a13_data;
wire [`DWIDTH-1:0] a14_data;
wire [`DWIDTH-1:0] a15_data;
wire [`DWIDTH-1:0] a16_data;
wire [`DWIDTH-1:0] a17_data;
wire [`DWIDTH-1:0] a18_data;
wire [`DWIDTH-1:0] a19_data;
wire [`DWIDTH-1:0] a20_data;
wire [`DWIDTH-1:0] a21_data;
wire [`DWIDTH-1:0] a22_data;
wire [`DWIDTH-1:0] a23_data;
wire [`DWIDTH-1:0] a24_data;
wire [`DWIDTH-1:0] a25_data;
wire [`DWIDTH-1:0] a26_data;
wire [`DWIDTH-1:0] a27_data;
wire [`DWIDTH-1:0] a28_data;
wire [`DWIDTH-1:0] a29_data;
wire [`DWIDTH-1:0] a30_data;
wire [`DWIDTH-1:0] a31_data;
wire [`DWIDTH-1:0] b0_data;
wire [`DWIDTH-1:0] b1_data;
wire [`DWIDTH-1:0] b2_data;
wire [`DWIDTH-1:0] b3_data;
wire [`DWIDTH-1:0] b4_data;
wire [`DWIDTH-1:0] b5_data;
wire [`DWIDTH-1:0] b6_data;
wire [`DWIDTH-1:0] b7_data;
wire [`DWIDTH-1:0] b8_data;
wire [`DWIDTH-1:0] b9_data;
wire [`DWIDTH-1:0] b10_data;
wire [`DWIDTH-1:0] b11_data;
wire [`DWIDTH-1:0] b12_data;
wire [`DWIDTH-1:0] b13_data;
wire [`DWIDTH-1:0] b14_data;
wire [`DWIDTH-1:0] b15_data;
wire [`DWIDTH-1:0] b16_data;
wire [`DWIDTH-1:0] b17_data;
wire [`DWIDTH-1:0] b18_data;
wire [`DWIDTH-1:0] b19_data;
wire [`DWIDTH-1:0] b20_data;
wire [`DWIDTH-1:0] b21_data;
wire [`DWIDTH-1:0] b22_data;
wire [`DWIDTH-1:0] b23_data;
wire [`DWIDTH-1:0] b24_data;
wire [`DWIDTH-1:0] b25_data;
wire [`DWIDTH-1:0] b26_data;
wire [`DWIDTH-1:0] b27_data;
wire [`DWIDTH-1:0] b28_data;
wire [`DWIDTH-1:0] b29_data;
wire [`DWIDTH-1:0] b30_data;
wire [`DWIDTH-1:0] b31_data;

//////////////////////////////////////////////////////////////////////////
// Logic to generate addresses to BRAM A
//////////////////////////////////////////////////////////////////////////
reg [`AWIDTH-1:0] a_addr;
reg a_mem_access; //flag that tells whether the matmul is trying to access memory or not

always @(posedge clk) begin
  //(clk_cnt >= a_loc*`MAT_MUL_SIZE+final_mat_mul_size) begin
  //Writing the line above to avoid multiplication:

  if (reset || ~start_mat_mul || (clk_cnt >= (a_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin
  
      a_addr <= address_mat_a-address_stride_a;
  
    a_mem_access <= 0;
  end
  //else if ((clk_cnt >= a_loc*`MAT_MUL_SIZE) && (clk_cnt < a_loc*`MAT_MUL_SIZE+final_mat_mul_size)) begin
  //Writing the line above to avoid multiplication:

  else if ((clk_cnt >= (a_loc<<`LOG2_MAT_MUL_SIZE)) && (clk_cnt < (a_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin
  
      a_addr <= a_addr + address_stride_a;
  
    a_mem_access <= 1;
  end
end

//////////////////////////////////////////////////////////////////////////
// Logic to generate valid signals for data coming from BRAM A
//////////////////////////////////////////////////////////////////////////
reg [7:0] a_mem_access_counter;
always @(posedge clk) begin
  if (reset || ~start_mat_mul) begin
    a_mem_access_counter <= 0;
  end
  else if (a_mem_access == 1) begin
    a_mem_access_counter <= a_mem_access_counter + 1;  
  end
  else begin
    a_mem_access_counter <= 0;
  end
end

wire a_data_valid; //flag that tells whether the data from memory is valid
assign a_data_valid = 
     ((validity_mask_a_cols_b_rows[0]==1'b0 && a_mem_access_counter==1) ||
      (validity_mask_a_cols_b_rows[1]==1'b0 && a_mem_access_counter==2) ||
      (validity_mask_a_cols_b_rows[2]==1'b0 && a_mem_access_counter==3) ||
      (validity_mask_a_cols_b_rows[3]==1'b0 && a_mem_access_counter==4) ||
      (validity_mask_a_cols_b_rows[4]==1'b0 && a_mem_access_counter==5) ||
      (validity_mask_a_cols_b_rows[5]==1'b0 && a_mem_access_counter==6) ||
      (validity_mask_a_cols_b_rows[6]==1'b0 && a_mem_access_counter==7) ||
      (validity_mask_a_cols_b_rows[7]==1'b0 && a_mem_access_counter==8) ||
      (validity_mask_a_cols_b_rows[8]==1'b0 && a_mem_access_counter==9) ||
      (validity_mask_a_cols_b_rows[9]==1'b0 && a_mem_access_counter==10) ||
      (validity_mask_a_cols_b_rows[10]==1'b0 && a_mem_access_counter==11) ||
      (validity_mask_a_cols_b_rows[11]==1'b0 && a_mem_access_counter==12) ||
      (validity_mask_a_cols_b_rows[12]==1'b0 && a_mem_access_counter==13) ||
      (validity_mask_a_cols_b_rows[13]==1'b0 && a_mem_access_counter==14) ||
      (validity_mask_a_cols_b_rows[14]==1'b0 && a_mem_access_counter==15) ||
      (validity_mask_a_cols_b_rows[15]==1'b0 && a_mem_access_counter==16) ||
      (validity_mask_a_cols_b_rows[16]==1'b0 && a_mem_access_counter==17) ||
      (validity_mask_a_cols_b_rows[17]==1'b0 && a_mem_access_counter==18) ||
      (validity_mask_a_cols_b_rows[18]==1'b0 && a_mem_access_counter==19) ||
      (validity_mask_a_cols_b_rows[19]==1'b0 && a_mem_access_counter==20) ||
      (validity_mask_a_cols_b_rows[20]==1'b0 && a_mem_access_counter==21) ||
      (validity_mask_a_cols_b_rows[21]==1'b0 && a_mem_access_counter==22) ||
      (validity_mask_a_cols_b_rows[22]==1'b0 && a_mem_access_counter==23) ||
      (validity_mask_a_cols_b_rows[23]==1'b0 && a_mem_access_counter==24) ||
      (validity_mask_a_cols_b_rows[24]==1'b0 && a_mem_access_counter==25) ||
      (validity_mask_a_cols_b_rows[25]==1'b0 && a_mem_access_counter==26) ||
      (validity_mask_a_cols_b_rows[26]==1'b0 && a_mem_access_counter==27) ||
      (validity_mask_a_cols_b_rows[27]==1'b0 && a_mem_access_counter==28) ||
      (validity_mask_a_cols_b_rows[28]==1'b0 && a_mem_access_counter==29) ||
      (validity_mask_a_cols_b_rows[29]==1'b0 && a_mem_access_counter==30) ||
      (validity_mask_a_cols_b_rows[30]==1'b0 && a_mem_access_counter==31) ||
      (validity_mask_a_cols_b_rows[31]==1'b0 && a_mem_access_counter==32)) ?
    
    1'b0 : (a_mem_access_counter >= `MEM_ACCESS_LATENCY);

//////////////////////////////////////////////////////////////////////////
// Logic to delay certain parts of the data received from BRAM A (systolic data setup)
//////////////////////////////////////////////////////////////////////////
assign a0_data = a_data[1*`DWIDTH-1:0*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[0]}};
assign a1_data = a_data[2*`DWIDTH-1:1*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[1]}};
assign a2_data = a_data[3*`DWIDTH-1:2*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[2]}};
assign a3_data = a_data[4*`DWIDTH-1:3*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[3]}};
assign a4_data = a_data[5*`DWIDTH-1:4*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[4]}};
assign a5_data = a_data[6*`DWIDTH-1:5*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[5]}};
assign a6_data = a_data[7*`DWIDTH-1:6*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[6]}};
assign a7_data = a_data[8*`DWIDTH-1:7*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[7]}};
assign a8_data = a_data[9*`DWIDTH-1:8*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[8]}};
assign a9_data = a_data[10*`DWIDTH-1:9*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[9]}};
assign a10_data = a_data[11*`DWIDTH-1:10*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[10]}};
assign a11_data = a_data[12*`DWIDTH-1:11*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[11]}};
assign a12_data = a_data[13*`DWIDTH-1:12*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[12]}};
assign a13_data = a_data[14*`DWIDTH-1:13*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[13]}};
assign a14_data = a_data[15*`DWIDTH-1:14*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[14]}};
assign a15_data = a_data[16*`DWIDTH-1:15*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[15]}};
assign a16_data = a_data[17*`DWIDTH-1:16*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[16]}};
assign a17_data = a_data[18*`DWIDTH-1:17*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[17]}};
assign a18_data = a_data[19*`DWIDTH-1:18*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[18]}};
assign a19_data = a_data[20*`DWIDTH-1:19*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[19]}};
assign a20_data = a_data[21*`DWIDTH-1:20*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[20]}};
assign a21_data = a_data[22*`DWIDTH-1:21*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[21]}};
assign a22_data = a_data[23*`DWIDTH-1:22*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[22]}};
assign a23_data = a_data[24*`DWIDTH-1:23*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[23]}};
assign a24_data = a_data[25*`DWIDTH-1:24*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[24]}};
assign a25_data = a_data[26*`DWIDTH-1:25*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[25]}};
assign a26_data = a_data[27*`DWIDTH-1:26*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[26]}};
assign a27_data = a_data[28*`DWIDTH-1:27*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[27]}};
assign a28_data = a_data[29*`DWIDTH-1:28*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[28]}};
assign a29_data = a_data[30*`DWIDTH-1:29*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[29]}};
assign a30_data = a_data[31*`DWIDTH-1:30*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[30]}};
assign a31_data = a_data[32*`DWIDTH-1:31*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[31]}};

reg [`DWIDTH-1:0] a1_data_delayed_1;
reg [`DWIDTH-1:0] a2_data_delayed_1;
reg [`DWIDTH-1:0] a2_data_delayed_2;
reg [`DWIDTH-1:0] a3_data_delayed_1;
reg [`DWIDTH-1:0] a3_data_delayed_2;
reg [`DWIDTH-1:0] a3_data_delayed_3;
reg [`DWIDTH-1:0] a4_data_delayed_1;
reg [`DWIDTH-1:0] a4_data_delayed_2;
reg [`DWIDTH-1:0] a4_data_delayed_3;
reg [`DWIDTH-1:0] a4_data_delayed_4;
reg [`DWIDTH-1:0] a5_data_delayed_1;
reg [`DWIDTH-1:0] a5_data_delayed_2;
reg [`DWIDTH-1:0] a5_data_delayed_3;
reg [`DWIDTH-1:0] a5_data_delayed_4;
reg [`DWIDTH-1:0] a5_data_delayed_5;
reg [`DWIDTH-1:0] a6_data_delayed_1;
reg [`DWIDTH-1:0] a6_data_delayed_2;
reg [`DWIDTH-1:0] a6_data_delayed_3;
reg [`DWIDTH-1:0] a6_data_delayed_4;
reg [`DWIDTH-1:0] a6_data_delayed_5;
reg [`DWIDTH-1:0] a6_data_delayed_6;
reg [`DWIDTH-1:0] a7_data_delayed_1;
reg [`DWIDTH-1:0] a7_data_delayed_2;
reg [`DWIDTH-1:0] a7_data_delayed_3;
reg [`DWIDTH-1:0] a7_data_delayed_4;
reg [`DWIDTH-1:0] a7_data_delayed_5;
reg [`DWIDTH-1:0] a7_data_delayed_6;
reg [`DWIDTH-1:0] a7_data_delayed_7;
reg [`DWIDTH-1:0] a8_data_delayed_1;
reg [`DWIDTH-1:0] a8_data_delayed_2;
reg [`DWIDTH-1:0] a8_data_delayed_3;
reg [`DWIDTH-1:0] a8_data_delayed_4;
reg [`DWIDTH-1:0] a8_data_delayed_5;
reg [`DWIDTH-1:0] a8_data_delayed_6;
reg [`DWIDTH-1:0] a8_data_delayed_7;
reg [`DWIDTH-1:0] a8_data_delayed_8;
reg [`DWIDTH-1:0] a9_data_delayed_1;
reg [`DWIDTH-1:0] a9_data_delayed_2;
reg [`DWIDTH-1:0] a9_data_delayed_3;
reg [`DWIDTH-1:0] a9_data_delayed_4;
reg [`DWIDTH-1:0] a9_data_delayed_5;
reg [`DWIDTH-1:0] a9_data_delayed_6;
reg [`DWIDTH-1:0] a9_data_delayed_7;
reg [`DWIDTH-1:0] a9_data_delayed_8;
reg [`DWIDTH-1:0] a9_data_delayed_9;
reg [`DWIDTH-1:0] a10_data_delayed_1;
reg [`DWIDTH-1:0] a10_data_delayed_2;
reg [`DWIDTH-1:0] a10_data_delayed_3;
reg [`DWIDTH-1:0] a10_data_delayed_4;
reg [`DWIDTH-1:0] a10_data_delayed_5;
reg [`DWIDTH-1:0] a10_data_delayed_6;
reg [`DWIDTH-1:0] a10_data_delayed_7;
reg [`DWIDTH-1:0] a10_data_delayed_8;
reg [`DWIDTH-1:0] a10_data_delayed_9;
reg [`DWIDTH-1:0] a10_data_delayed_10;
reg [`DWIDTH-1:0] a11_data_delayed_1;
reg [`DWIDTH-1:0] a11_data_delayed_2;
reg [`DWIDTH-1:0] a11_data_delayed_3;
reg [`DWIDTH-1:0] a11_data_delayed_4;
reg [`DWIDTH-1:0] a11_data_delayed_5;
reg [`DWIDTH-1:0] a11_data_delayed_6;
reg [`DWIDTH-1:0] a11_data_delayed_7;
reg [`DWIDTH-1:0] a11_data_delayed_8;
reg [`DWIDTH-1:0] a11_data_delayed_9;
reg [`DWIDTH-1:0] a11_data_delayed_10;
reg [`DWIDTH-1:0] a11_data_delayed_11;
reg [`DWIDTH-1:0] a12_data_delayed_1;
reg [`DWIDTH-1:0] a12_data_delayed_2;
reg [`DWIDTH-1:0] a12_data_delayed_3;
reg [`DWIDTH-1:0] a12_data_delayed_4;
reg [`DWIDTH-1:0] a12_data_delayed_5;
reg [`DWIDTH-1:0] a12_data_delayed_6;
reg [`DWIDTH-1:0] a12_data_delayed_7;
reg [`DWIDTH-1:0] a12_data_delayed_8;
reg [`DWIDTH-1:0] a12_data_delayed_9;
reg [`DWIDTH-1:0] a12_data_delayed_10;
reg [`DWIDTH-1:0] a12_data_delayed_11;
reg [`DWIDTH-1:0] a12_data_delayed_12;
reg [`DWIDTH-1:0] a13_data_delayed_1;
reg [`DWIDTH-1:0] a13_data_delayed_2;
reg [`DWIDTH-1:0] a13_data_delayed_3;
reg [`DWIDTH-1:0] a13_data_delayed_4;
reg [`DWIDTH-1:0] a13_data_delayed_5;
reg [`DWIDTH-1:0] a13_data_delayed_6;
reg [`DWIDTH-1:0] a13_data_delayed_7;
reg [`DWIDTH-1:0] a13_data_delayed_8;
reg [`DWIDTH-1:0] a13_data_delayed_9;
reg [`DWIDTH-1:0] a13_data_delayed_10;
reg [`DWIDTH-1:0] a13_data_delayed_11;
reg [`DWIDTH-1:0] a13_data_delayed_12;
reg [`DWIDTH-1:0] a13_data_delayed_13;
reg [`DWIDTH-1:0] a14_data_delayed_1;
reg [`DWIDTH-1:0] a14_data_delayed_2;
reg [`DWIDTH-1:0] a14_data_delayed_3;
reg [`DWIDTH-1:0] a14_data_delayed_4;
reg [`DWIDTH-1:0] a14_data_delayed_5;
reg [`DWIDTH-1:0] a14_data_delayed_6;
reg [`DWIDTH-1:0] a14_data_delayed_7;
reg [`DWIDTH-1:0] a14_data_delayed_8;
reg [`DWIDTH-1:0] a14_data_delayed_9;
reg [`DWIDTH-1:0] a14_data_delayed_10;
reg [`DWIDTH-1:0] a14_data_delayed_11;
reg [`DWIDTH-1:0] a14_data_delayed_12;
reg [`DWIDTH-1:0] a14_data_delayed_13;
reg [`DWIDTH-1:0] a14_data_delayed_14;
reg [`DWIDTH-1:0] a15_data_delayed_1;
reg [`DWIDTH-1:0] a15_data_delayed_2;
reg [`DWIDTH-1:0] a15_data_delayed_3;
reg [`DWIDTH-1:0] a15_data_delayed_4;
reg [`DWIDTH-1:0] a15_data_delayed_5;
reg [`DWIDTH-1:0] a15_data_delayed_6;
reg [`DWIDTH-1:0] a15_data_delayed_7;
reg [`DWIDTH-1:0] a15_data_delayed_8;
reg [`DWIDTH-1:0] a15_data_delayed_9;
reg [`DWIDTH-1:0] a15_data_delayed_10;
reg [`DWIDTH-1:0] a15_data_delayed_11;
reg [`DWIDTH-1:0] a15_data_delayed_12;
reg [`DWIDTH-1:0] a15_data_delayed_13;
reg [`DWIDTH-1:0] a15_data_delayed_14;
reg [`DWIDTH-1:0] a15_data_delayed_15;
reg [`DWIDTH-1:0] a16_data_delayed_1;
reg [`DWIDTH-1:0] a16_data_delayed_2;
reg [`DWIDTH-1:0] a16_data_delayed_3;
reg [`DWIDTH-1:0] a16_data_delayed_4;
reg [`DWIDTH-1:0] a16_data_delayed_5;
reg [`DWIDTH-1:0] a16_data_delayed_6;
reg [`DWIDTH-1:0] a16_data_delayed_7;
reg [`DWIDTH-1:0] a16_data_delayed_8;
reg [`DWIDTH-1:0] a16_data_delayed_9;
reg [`DWIDTH-1:0] a16_data_delayed_10;
reg [`DWIDTH-1:0] a16_data_delayed_11;
reg [`DWIDTH-1:0] a16_data_delayed_12;
reg [`DWIDTH-1:0] a16_data_delayed_13;
reg [`DWIDTH-1:0] a16_data_delayed_14;
reg [`DWIDTH-1:0] a16_data_delayed_15;
reg [`DWIDTH-1:0] a16_data_delayed_16;
reg [`DWIDTH-1:0] a17_data_delayed_1;
reg [`DWIDTH-1:0] a17_data_delayed_2;
reg [`DWIDTH-1:0] a17_data_delayed_3;
reg [`DWIDTH-1:0] a17_data_delayed_4;
reg [`DWIDTH-1:0] a17_data_delayed_5;
reg [`DWIDTH-1:0] a17_data_delayed_6;
reg [`DWIDTH-1:0] a17_data_delayed_7;
reg [`DWIDTH-1:0] a17_data_delayed_8;
reg [`DWIDTH-1:0] a17_data_delayed_9;
reg [`DWIDTH-1:0] a17_data_delayed_10;
reg [`DWIDTH-1:0] a17_data_delayed_11;
reg [`DWIDTH-1:0] a17_data_delayed_12;
reg [`DWIDTH-1:0] a17_data_delayed_13;
reg [`DWIDTH-1:0] a17_data_delayed_14;
reg [`DWIDTH-1:0] a17_data_delayed_15;
reg [`DWIDTH-1:0] a17_data_delayed_16;
reg [`DWIDTH-1:0] a17_data_delayed_17;
reg [`DWIDTH-1:0] a18_data_delayed_1;
reg [`DWIDTH-1:0] a18_data_delayed_2;
reg [`DWIDTH-1:0] a18_data_delayed_3;
reg [`DWIDTH-1:0] a18_data_delayed_4;
reg [`DWIDTH-1:0] a18_data_delayed_5;
reg [`DWIDTH-1:0] a18_data_delayed_6;
reg [`DWIDTH-1:0] a18_data_delayed_7;
reg [`DWIDTH-1:0] a18_data_delayed_8;
reg [`DWIDTH-1:0] a18_data_delayed_9;
reg [`DWIDTH-1:0] a18_data_delayed_10;
reg [`DWIDTH-1:0] a18_data_delayed_11;
reg [`DWIDTH-1:0] a18_data_delayed_12;
reg [`DWIDTH-1:0] a18_data_delayed_13;
reg [`DWIDTH-1:0] a18_data_delayed_14;
reg [`DWIDTH-1:0] a18_data_delayed_15;
reg [`DWIDTH-1:0] a18_data_delayed_16;
reg [`DWIDTH-1:0] a18_data_delayed_17;
reg [`DWIDTH-1:0] a18_data_delayed_18;
reg [`DWIDTH-1:0] a19_data_delayed_1;
reg [`DWIDTH-1:0] a19_data_delayed_2;
reg [`DWIDTH-1:0] a19_data_delayed_3;
reg [`DWIDTH-1:0] a19_data_delayed_4;
reg [`DWIDTH-1:0] a19_data_delayed_5;
reg [`DWIDTH-1:0] a19_data_delayed_6;
reg [`DWIDTH-1:0] a19_data_delayed_7;
reg [`DWIDTH-1:0] a19_data_delayed_8;
reg [`DWIDTH-1:0] a19_data_delayed_9;
reg [`DWIDTH-1:0] a19_data_delayed_10;
reg [`DWIDTH-1:0] a19_data_delayed_11;
reg [`DWIDTH-1:0] a19_data_delayed_12;
reg [`DWIDTH-1:0] a19_data_delayed_13;
reg [`DWIDTH-1:0] a19_data_delayed_14;
reg [`DWIDTH-1:0] a19_data_delayed_15;
reg [`DWIDTH-1:0] a19_data_delayed_16;
reg [`DWIDTH-1:0] a19_data_delayed_17;
reg [`DWIDTH-1:0] a19_data_delayed_18;
reg [`DWIDTH-1:0] a19_data_delayed_19;
reg [`DWIDTH-1:0] a20_data_delayed_1;
reg [`DWIDTH-1:0] a20_data_delayed_2;
reg [`DWIDTH-1:0] a20_data_delayed_3;
reg [`DWIDTH-1:0] a20_data_delayed_4;
reg [`DWIDTH-1:0] a20_data_delayed_5;
reg [`DWIDTH-1:0] a20_data_delayed_6;
reg [`DWIDTH-1:0] a20_data_delayed_7;
reg [`DWIDTH-1:0] a20_data_delayed_8;
reg [`DWIDTH-1:0] a20_data_delayed_9;
reg [`DWIDTH-1:0] a20_data_delayed_10;
reg [`DWIDTH-1:0] a20_data_delayed_11;
reg [`DWIDTH-1:0] a20_data_delayed_12;
reg [`DWIDTH-1:0] a20_data_delayed_13;
reg [`DWIDTH-1:0] a20_data_delayed_14;
reg [`DWIDTH-1:0] a20_data_delayed_15;
reg [`DWIDTH-1:0] a20_data_delayed_16;
reg [`DWIDTH-1:0] a20_data_delayed_17;
reg [`DWIDTH-1:0] a20_data_delayed_18;
reg [`DWIDTH-1:0] a20_data_delayed_19;
reg [`DWIDTH-1:0] a20_data_delayed_20;
reg [`DWIDTH-1:0] a21_data_delayed_1;
reg [`DWIDTH-1:0] a21_data_delayed_2;
reg [`DWIDTH-1:0] a21_data_delayed_3;
reg [`DWIDTH-1:0] a21_data_delayed_4;
reg [`DWIDTH-1:0] a21_data_delayed_5;
reg [`DWIDTH-1:0] a21_data_delayed_6;
reg [`DWIDTH-1:0] a21_data_delayed_7;
reg [`DWIDTH-1:0] a21_data_delayed_8;
reg [`DWIDTH-1:0] a21_data_delayed_9;
reg [`DWIDTH-1:0] a21_data_delayed_10;
reg [`DWIDTH-1:0] a21_data_delayed_11;
reg [`DWIDTH-1:0] a21_data_delayed_12;
reg [`DWIDTH-1:0] a21_data_delayed_13;
reg [`DWIDTH-1:0] a21_data_delayed_14;
reg [`DWIDTH-1:0] a21_data_delayed_15;
reg [`DWIDTH-1:0] a21_data_delayed_16;
reg [`DWIDTH-1:0] a21_data_delayed_17;
reg [`DWIDTH-1:0] a21_data_delayed_18;
reg [`DWIDTH-1:0] a21_data_delayed_19;
reg [`DWIDTH-1:0] a21_data_delayed_20;
reg [`DWIDTH-1:0] a21_data_delayed_21;
reg [`DWIDTH-1:0] a22_data_delayed_1;
reg [`DWIDTH-1:0] a22_data_delayed_2;
reg [`DWIDTH-1:0] a22_data_delayed_3;
reg [`DWIDTH-1:0] a22_data_delayed_4;
reg [`DWIDTH-1:0] a22_data_delayed_5;
reg [`DWIDTH-1:0] a22_data_delayed_6;
reg [`DWIDTH-1:0] a22_data_delayed_7;
reg [`DWIDTH-1:0] a22_data_delayed_8;
reg [`DWIDTH-1:0] a22_data_delayed_9;
reg [`DWIDTH-1:0] a22_data_delayed_10;
reg [`DWIDTH-1:0] a22_data_delayed_11;
reg [`DWIDTH-1:0] a22_data_delayed_12;
reg [`DWIDTH-1:0] a22_data_delayed_13;
reg [`DWIDTH-1:0] a22_data_delayed_14;
reg [`DWIDTH-1:0] a22_data_delayed_15;
reg [`DWIDTH-1:0] a22_data_delayed_16;
reg [`DWIDTH-1:0] a22_data_delayed_17;
reg [`DWIDTH-1:0] a22_data_delayed_18;
reg [`DWIDTH-1:0] a22_data_delayed_19;
reg [`DWIDTH-1:0] a22_data_delayed_20;
reg [`DWIDTH-1:0] a22_data_delayed_21;
reg [`DWIDTH-1:0] a22_data_delayed_22;
reg [`DWIDTH-1:0] a23_data_delayed_1;
reg [`DWIDTH-1:0] a23_data_delayed_2;
reg [`DWIDTH-1:0] a23_data_delayed_3;
reg [`DWIDTH-1:0] a23_data_delayed_4;
reg [`DWIDTH-1:0] a23_data_delayed_5;
reg [`DWIDTH-1:0] a23_data_delayed_6;
reg [`DWIDTH-1:0] a23_data_delayed_7;
reg [`DWIDTH-1:0] a23_data_delayed_8;
reg [`DWIDTH-1:0] a23_data_delayed_9;
reg [`DWIDTH-1:0] a23_data_delayed_10;
reg [`DWIDTH-1:0] a23_data_delayed_11;
reg [`DWIDTH-1:0] a23_data_delayed_12;
reg [`DWIDTH-1:0] a23_data_delayed_13;
reg [`DWIDTH-1:0] a23_data_delayed_14;
reg [`DWIDTH-1:0] a23_data_delayed_15;
reg [`DWIDTH-1:0] a23_data_delayed_16;
reg [`DWIDTH-1:0] a23_data_delayed_17;
reg [`DWIDTH-1:0] a23_data_delayed_18;
reg [`DWIDTH-1:0] a23_data_delayed_19;
reg [`DWIDTH-1:0] a23_data_delayed_20;
reg [`DWIDTH-1:0] a23_data_delayed_21;
reg [`DWIDTH-1:0] a23_data_delayed_22;
reg [`DWIDTH-1:0] a23_data_delayed_23;
reg [`DWIDTH-1:0] a24_data_delayed_1;
reg [`DWIDTH-1:0] a24_data_delayed_2;
reg [`DWIDTH-1:0] a24_data_delayed_3;
reg [`DWIDTH-1:0] a24_data_delayed_4;
reg [`DWIDTH-1:0] a24_data_delayed_5;
reg [`DWIDTH-1:0] a24_data_delayed_6;
reg [`DWIDTH-1:0] a24_data_delayed_7;
reg [`DWIDTH-1:0] a24_data_delayed_8;
reg [`DWIDTH-1:0] a24_data_delayed_9;
reg [`DWIDTH-1:0] a24_data_delayed_10;
reg [`DWIDTH-1:0] a24_data_delayed_11;
reg [`DWIDTH-1:0] a24_data_delayed_12;
reg [`DWIDTH-1:0] a24_data_delayed_13;
reg [`DWIDTH-1:0] a24_data_delayed_14;
reg [`DWIDTH-1:0] a24_data_delayed_15;
reg [`DWIDTH-1:0] a24_data_delayed_16;
reg [`DWIDTH-1:0] a24_data_delayed_17;
reg [`DWIDTH-1:0] a24_data_delayed_18;
reg [`DWIDTH-1:0] a24_data_delayed_19;
reg [`DWIDTH-1:0] a24_data_delayed_20;
reg [`DWIDTH-1:0] a24_data_delayed_21;
reg [`DWIDTH-1:0] a24_data_delayed_22;
reg [`DWIDTH-1:0] a24_data_delayed_23;
reg [`DWIDTH-1:0] a24_data_delayed_24;
reg [`DWIDTH-1:0] a25_data_delayed_1;
reg [`DWIDTH-1:0] a25_data_delayed_2;
reg [`DWIDTH-1:0] a25_data_delayed_3;
reg [`DWIDTH-1:0] a25_data_delayed_4;
reg [`DWIDTH-1:0] a25_data_delayed_5;
reg [`DWIDTH-1:0] a25_data_delayed_6;
reg [`DWIDTH-1:0] a25_data_delayed_7;
reg [`DWIDTH-1:0] a25_data_delayed_8;
reg [`DWIDTH-1:0] a25_data_delayed_9;
reg [`DWIDTH-1:0] a25_data_delayed_10;
reg [`DWIDTH-1:0] a25_data_delayed_11;
reg [`DWIDTH-1:0] a25_data_delayed_12;
reg [`DWIDTH-1:0] a25_data_delayed_13;
reg [`DWIDTH-1:0] a25_data_delayed_14;
reg [`DWIDTH-1:0] a25_data_delayed_15;
reg [`DWIDTH-1:0] a25_data_delayed_16;
reg [`DWIDTH-1:0] a25_data_delayed_17;
reg [`DWIDTH-1:0] a25_data_delayed_18;
reg [`DWIDTH-1:0] a25_data_delayed_19;
reg [`DWIDTH-1:0] a25_data_delayed_20;
reg [`DWIDTH-1:0] a25_data_delayed_21;
reg [`DWIDTH-1:0] a25_data_delayed_22;
reg [`DWIDTH-1:0] a25_data_delayed_23;
reg [`DWIDTH-1:0] a25_data_delayed_24;
reg [`DWIDTH-1:0] a25_data_delayed_25;
reg [`DWIDTH-1:0] a26_data_delayed_1;
reg [`DWIDTH-1:0] a26_data_delayed_2;
reg [`DWIDTH-1:0] a26_data_delayed_3;
reg [`DWIDTH-1:0] a26_data_delayed_4;
reg [`DWIDTH-1:0] a26_data_delayed_5;
reg [`DWIDTH-1:0] a26_data_delayed_6;
reg [`DWIDTH-1:0] a26_data_delayed_7;
reg [`DWIDTH-1:0] a26_data_delayed_8;
reg [`DWIDTH-1:0] a26_data_delayed_9;
reg [`DWIDTH-1:0] a26_data_delayed_10;
reg [`DWIDTH-1:0] a26_data_delayed_11;
reg [`DWIDTH-1:0] a26_data_delayed_12;
reg [`DWIDTH-1:0] a26_data_delayed_13;
reg [`DWIDTH-1:0] a26_data_delayed_14;
reg [`DWIDTH-1:0] a26_data_delayed_15;
reg [`DWIDTH-1:0] a26_data_delayed_16;
reg [`DWIDTH-1:0] a26_data_delayed_17;
reg [`DWIDTH-1:0] a26_data_delayed_18;
reg [`DWIDTH-1:0] a26_data_delayed_19;
reg [`DWIDTH-1:0] a26_data_delayed_20;
reg [`DWIDTH-1:0] a26_data_delayed_21;
reg [`DWIDTH-1:0] a26_data_delayed_22;
reg [`DWIDTH-1:0] a26_data_delayed_23;
reg [`DWIDTH-1:0] a26_data_delayed_24;
reg [`DWIDTH-1:0] a26_data_delayed_25;
reg [`DWIDTH-1:0] a26_data_delayed_26;
reg [`DWIDTH-1:0] a27_data_delayed_1;
reg [`DWIDTH-1:0] a27_data_delayed_2;
reg [`DWIDTH-1:0] a27_data_delayed_3;
reg [`DWIDTH-1:0] a27_data_delayed_4;
reg [`DWIDTH-1:0] a27_data_delayed_5;
reg [`DWIDTH-1:0] a27_data_delayed_6;
reg [`DWIDTH-1:0] a27_data_delayed_7;
reg [`DWIDTH-1:0] a27_data_delayed_8;
reg [`DWIDTH-1:0] a27_data_delayed_9;
reg [`DWIDTH-1:0] a27_data_delayed_10;
reg [`DWIDTH-1:0] a27_data_delayed_11;
reg [`DWIDTH-1:0] a27_data_delayed_12;
reg [`DWIDTH-1:0] a27_data_delayed_13;
reg [`DWIDTH-1:0] a27_data_delayed_14;
reg [`DWIDTH-1:0] a27_data_delayed_15;
reg [`DWIDTH-1:0] a27_data_delayed_16;
reg [`DWIDTH-1:0] a27_data_delayed_17;
reg [`DWIDTH-1:0] a27_data_delayed_18;
reg [`DWIDTH-1:0] a27_data_delayed_19;
reg [`DWIDTH-1:0] a27_data_delayed_20;
reg [`DWIDTH-1:0] a27_data_delayed_21;
reg [`DWIDTH-1:0] a27_data_delayed_22;
reg [`DWIDTH-1:0] a27_data_delayed_23;
reg [`DWIDTH-1:0] a27_data_delayed_24;
reg [`DWIDTH-1:0] a27_data_delayed_25;
reg [`DWIDTH-1:0] a27_data_delayed_26;
reg [`DWIDTH-1:0] a27_data_delayed_27;
reg [`DWIDTH-1:0] a28_data_delayed_1;
reg [`DWIDTH-1:0] a28_data_delayed_2;
reg [`DWIDTH-1:0] a28_data_delayed_3;
reg [`DWIDTH-1:0] a28_data_delayed_4;
reg [`DWIDTH-1:0] a28_data_delayed_5;
reg [`DWIDTH-1:0] a28_data_delayed_6;
reg [`DWIDTH-1:0] a28_data_delayed_7;
reg [`DWIDTH-1:0] a28_data_delayed_8;
reg [`DWIDTH-1:0] a28_data_delayed_9;
reg [`DWIDTH-1:0] a28_data_delayed_10;
reg [`DWIDTH-1:0] a28_data_delayed_11;
reg [`DWIDTH-1:0] a28_data_delayed_12;
reg [`DWIDTH-1:0] a28_data_delayed_13;
reg [`DWIDTH-1:0] a28_data_delayed_14;
reg [`DWIDTH-1:0] a28_data_delayed_15;
reg [`DWIDTH-1:0] a28_data_delayed_16;
reg [`DWIDTH-1:0] a28_data_delayed_17;
reg [`DWIDTH-1:0] a28_data_delayed_18;
reg [`DWIDTH-1:0] a28_data_delayed_19;
reg [`DWIDTH-1:0] a28_data_delayed_20;
reg [`DWIDTH-1:0] a28_data_delayed_21;
reg [`DWIDTH-1:0] a28_data_delayed_22;
reg [`DWIDTH-1:0] a28_data_delayed_23;
reg [`DWIDTH-1:0] a28_data_delayed_24;
reg [`DWIDTH-1:0] a28_data_delayed_25;
reg [`DWIDTH-1:0] a28_data_delayed_26;
reg [`DWIDTH-1:0] a28_data_delayed_27;
reg [`DWIDTH-1:0] a28_data_delayed_28;
reg [`DWIDTH-1:0] a29_data_delayed_1;
reg [`DWIDTH-1:0] a29_data_delayed_2;
reg [`DWIDTH-1:0] a29_data_delayed_3;
reg [`DWIDTH-1:0] a29_data_delayed_4;
reg [`DWIDTH-1:0] a29_data_delayed_5;
reg [`DWIDTH-1:0] a29_data_delayed_6;
reg [`DWIDTH-1:0] a29_data_delayed_7;
reg [`DWIDTH-1:0] a29_data_delayed_8;
reg [`DWIDTH-1:0] a29_data_delayed_9;
reg [`DWIDTH-1:0] a29_data_delayed_10;
reg [`DWIDTH-1:0] a29_data_delayed_11;
reg [`DWIDTH-1:0] a29_data_delayed_12;
reg [`DWIDTH-1:0] a29_data_delayed_13;
reg [`DWIDTH-1:0] a29_data_delayed_14;
reg [`DWIDTH-1:0] a29_data_delayed_15;
reg [`DWIDTH-1:0] a29_data_delayed_16;
reg [`DWIDTH-1:0] a29_data_delayed_17;
reg [`DWIDTH-1:0] a29_data_delayed_18;
reg [`DWIDTH-1:0] a29_data_delayed_19;
reg [`DWIDTH-1:0] a29_data_delayed_20;
reg [`DWIDTH-1:0] a29_data_delayed_21;
reg [`DWIDTH-1:0] a29_data_delayed_22;
reg [`DWIDTH-1:0] a29_data_delayed_23;
reg [`DWIDTH-1:0] a29_data_delayed_24;
reg [`DWIDTH-1:0] a29_data_delayed_25;
reg [`DWIDTH-1:0] a29_data_delayed_26;
reg [`DWIDTH-1:0] a29_data_delayed_27;
reg [`DWIDTH-1:0] a29_data_delayed_28;
reg [`DWIDTH-1:0] a29_data_delayed_29;
reg [`DWIDTH-1:0] a30_data_delayed_1;
reg [`DWIDTH-1:0] a30_data_delayed_2;
reg [`DWIDTH-1:0] a30_data_delayed_3;
reg [`DWIDTH-1:0] a30_data_delayed_4;
reg [`DWIDTH-1:0] a30_data_delayed_5;
reg [`DWIDTH-1:0] a30_data_delayed_6;
reg [`DWIDTH-1:0] a30_data_delayed_7;
reg [`DWIDTH-1:0] a30_data_delayed_8;
reg [`DWIDTH-1:0] a30_data_delayed_9;
reg [`DWIDTH-1:0] a30_data_delayed_10;
reg [`DWIDTH-1:0] a30_data_delayed_11;
reg [`DWIDTH-1:0] a30_data_delayed_12;
reg [`DWIDTH-1:0] a30_data_delayed_13;
reg [`DWIDTH-1:0] a30_data_delayed_14;
reg [`DWIDTH-1:0] a30_data_delayed_15;
reg [`DWIDTH-1:0] a30_data_delayed_16;
reg [`DWIDTH-1:0] a30_data_delayed_17;
reg [`DWIDTH-1:0] a30_data_delayed_18;
reg [`DWIDTH-1:0] a30_data_delayed_19;
reg [`DWIDTH-1:0] a30_data_delayed_20;
reg [`DWIDTH-1:0] a30_data_delayed_21;
reg [`DWIDTH-1:0] a30_data_delayed_22;
reg [`DWIDTH-1:0] a30_data_delayed_23;
reg [`DWIDTH-1:0] a30_data_delayed_24;
reg [`DWIDTH-1:0] a30_data_delayed_25;
reg [`DWIDTH-1:0] a30_data_delayed_26;
reg [`DWIDTH-1:0] a30_data_delayed_27;
reg [`DWIDTH-1:0] a30_data_delayed_28;
reg [`DWIDTH-1:0] a30_data_delayed_29;
reg [`DWIDTH-1:0] a30_data_delayed_30;
reg [`DWIDTH-1:0] a31_data_delayed_1;
reg [`DWIDTH-1:0] a31_data_delayed_2;
reg [`DWIDTH-1:0] a31_data_delayed_3;
reg [`DWIDTH-1:0] a31_data_delayed_4;
reg [`DWIDTH-1:0] a31_data_delayed_5;
reg [`DWIDTH-1:0] a31_data_delayed_6;
reg [`DWIDTH-1:0] a31_data_delayed_7;
reg [`DWIDTH-1:0] a31_data_delayed_8;
reg [`DWIDTH-1:0] a31_data_delayed_9;
reg [`DWIDTH-1:0] a31_data_delayed_10;
reg [`DWIDTH-1:0] a31_data_delayed_11;
reg [`DWIDTH-1:0] a31_data_delayed_12;
reg [`DWIDTH-1:0] a31_data_delayed_13;
reg [`DWIDTH-1:0] a31_data_delayed_14;
reg [`DWIDTH-1:0] a31_data_delayed_15;
reg [`DWIDTH-1:0] a31_data_delayed_16;
reg [`DWIDTH-1:0] a31_data_delayed_17;
reg [`DWIDTH-1:0] a31_data_delayed_18;
reg [`DWIDTH-1:0] a31_data_delayed_19;
reg [`DWIDTH-1:0] a31_data_delayed_20;
reg [`DWIDTH-1:0] a31_data_delayed_21;
reg [`DWIDTH-1:0] a31_data_delayed_22;
reg [`DWIDTH-1:0] a31_data_delayed_23;
reg [`DWIDTH-1:0] a31_data_delayed_24;
reg [`DWIDTH-1:0] a31_data_delayed_25;
reg [`DWIDTH-1:0] a31_data_delayed_26;
reg [`DWIDTH-1:0] a31_data_delayed_27;
reg [`DWIDTH-1:0] a31_data_delayed_28;
reg [`DWIDTH-1:0] a31_data_delayed_29;
reg [`DWIDTH-1:0] a31_data_delayed_30;
reg [`DWIDTH-1:0] a31_data_delayed_31;


always @(posedge clk) begin
  if (reset || ~start_mat_mul || clk_cnt==0) begin
    a1_data_delayed_1 <= 0;
    a2_data_delayed_1 <= 0;
    a2_data_delayed_2 <= 0;
    a3_data_delayed_1 <= 0;
    a3_data_delayed_2 <= 0;
    a3_data_delayed_3 <= 0;
    a4_data_delayed_1 <= 0;
    a4_data_delayed_2 <= 0;
    a4_data_delayed_3 <= 0;
    a4_data_delayed_4 <= 0;
    a5_data_delayed_1 <= 0;
    a5_data_delayed_2 <= 0;
    a5_data_delayed_3 <= 0;
    a5_data_delayed_4 <= 0;
    a5_data_delayed_5 <= 0;
    a6_data_delayed_1 <= 0;
    a6_data_delayed_2 <= 0;
    a6_data_delayed_3 <= 0;
    a6_data_delayed_4 <= 0;
    a6_data_delayed_5 <= 0;
    a6_data_delayed_6 <= 0;
    a7_data_delayed_1 <= 0;
    a7_data_delayed_2 <= 0;
    a7_data_delayed_3 <= 0;
    a7_data_delayed_4 <= 0;
    a7_data_delayed_5 <= 0;
    a7_data_delayed_6 <= 0;
    a7_data_delayed_7 <= 0;
    a8_data_delayed_1 <= 0;
    a8_data_delayed_2 <= 0;
    a8_data_delayed_3 <= 0;
    a8_data_delayed_4 <= 0;
    a8_data_delayed_5 <= 0;
    a8_data_delayed_6 <= 0;
    a8_data_delayed_7 <= 0;
    a8_data_delayed_8 <= 0;
    a9_data_delayed_1 <= 0;
    a9_data_delayed_2 <= 0;
    a9_data_delayed_3 <= 0;
    a9_data_delayed_4 <= 0;
    a9_data_delayed_5 <= 0;
    a9_data_delayed_6 <= 0;
    a9_data_delayed_7 <= 0;
    a9_data_delayed_8 <= 0;
    a9_data_delayed_9 <= 0;
    a10_data_delayed_1 <= 0;
    a10_data_delayed_2 <= 0;
    a10_data_delayed_3 <= 0;
    a10_data_delayed_4 <= 0;
    a10_data_delayed_5 <= 0;
    a10_data_delayed_6 <= 0;
    a10_data_delayed_7 <= 0;
    a10_data_delayed_8 <= 0;
    a10_data_delayed_9 <= 0;
    a10_data_delayed_10 <= 0;
    a11_data_delayed_1 <= 0;
    a11_data_delayed_2 <= 0;
    a11_data_delayed_3 <= 0;
    a11_data_delayed_4 <= 0;
    a11_data_delayed_5 <= 0;
    a11_data_delayed_6 <= 0;
    a11_data_delayed_7 <= 0;
    a11_data_delayed_8 <= 0;
    a11_data_delayed_9 <= 0;
    a11_data_delayed_10 <= 0;
    a11_data_delayed_11 <= 0;
    a12_data_delayed_1 <= 0;
    a12_data_delayed_2 <= 0;
    a12_data_delayed_3 <= 0;
    a12_data_delayed_4 <= 0;
    a12_data_delayed_5 <= 0;
    a12_data_delayed_6 <= 0;
    a12_data_delayed_7 <= 0;
    a12_data_delayed_8 <= 0;
    a12_data_delayed_9 <= 0;
    a12_data_delayed_10 <= 0;
    a12_data_delayed_11 <= 0;
    a12_data_delayed_12 <= 0;
    a13_data_delayed_1 <= 0;
    a13_data_delayed_2 <= 0;
    a13_data_delayed_3 <= 0;
    a13_data_delayed_4 <= 0;
    a13_data_delayed_5 <= 0;
    a13_data_delayed_6 <= 0;
    a13_data_delayed_7 <= 0;
    a13_data_delayed_8 <= 0;
    a13_data_delayed_9 <= 0;
    a13_data_delayed_10 <= 0;
    a13_data_delayed_11 <= 0;
    a13_data_delayed_12 <= 0;
    a13_data_delayed_13 <= 0;
    a14_data_delayed_1 <= 0;
    a14_data_delayed_2 <= 0;
    a14_data_delayed_3 <= 0;
    a14_data_delayed_4 <= 0;
    a14_data_delayed_5 <= 0;
    a14_data_delayed_6 <= 0;
    a14_data_delayed_7 <= 0;
    a14_data_delayed_8 <= 0;
    a14_data_delayed_9 <= 0;
    a14_data_delayed_10 <= 0;
    a14_data_delayed_11 <= 0;
    a14_data_delayed_12 <= 0;
    a14_data_delayed_13 <= 0;
    a14_data_delayed_14 <= 0;
    a15_data_delayed_1 <= 0;
    a15_data_delayed_2 <= 0;
    a15_data_delayed_3 <= 0;
    a15_data_delayed_4 <= 0;
    a15_data_delayed_5 <= 0;
    a15_data_delayed_6 <= 0;
    a15_data_delayed_7 <= 0;
    a15_data_delayed_8 <= 0;
    a15_data_delayed_9 <= 0;
    a15_data_delayed_10 <= 0;
    a15_data_delayed_11 <= 0;
    a15_data_delayed_12 <= 0;
    a15_data_delayed_13 <= 0;
    a15_data_delayed_14 <= 0;
    a15_data_delayed_15 <= 0;
    a16_data_delayed_1 <= 0;
    a16_data_delayed_2 <= 0;
    a16_data_delayed_3 <= 0;
    a16_data_delayed_4 <= 0;
    a16_data_delayed_5 <= 0;
    a16_data_delayed_6 <= 0;
    a16_data_delayed_7 <= 0;
    a16_data_delayed_8 <= 0;
    a16_data_delayed_9 <= 0;
    a16_data_delayed_10 <= 0;
    a16_data_delayed_11 <= 0;
    a16_data_delayed_12 <= 0;
    a16_data_delayed_13 <= 0;
    a16_data_delayed_14 <= 0;
    a16_data_delayed_15 <= 0;
    a16_data_delayed_16 <= 0;
    a17_data_delayed_1 <= 0;
    a17_data_delayed_2 <= 0;
    a17_data_delayed_3 <= 0;
    a17_data_delayed_4 <= 0;
    a17_data_delayed_5 <= 0;
    a17_data_delayed_6 <= 0;
    a17_data_delayed_7 <= 0;
    a17_data_delayed_8 <= 0;
    a17_data_delayed_9 <= 0;
    a17_data_delayed_10 <= 0;
    a17_data_delayed_11 <= 0;
    a17_data_delayed_12 <= 0;
    a17_data_delayed_13 <= 0;
    a17_data_delayed_14 <= 0;
    a17_data_delayed_15 <= 0;
    a17_data_delayed_16 <= 0;
    a17_data_delayed_17 <= 0;
    a18_data_delayed_1 <= 0;
    a18_data_delayed_2 <= 0;
    a18_data_delayed_3 <= 0;
    a18_data_delayed_4 <= 0;
    a18_data_delayed_5 <= 0;
    a18_data_delayed_6 <= 0;
    a18_data_delayed_7 <= 0;
    a18_data_delayed_8 <= 0;
    a18_data_delayed_9 <= 0;
    a18_data_delayed_10 <= 0;
    a18_data_delayed_11 <= 0;
    a18_data_delayed_12 <= 0;
    a18_data_delayed_13 <= 0;
    a18_data_delayed_14 <= 0;
    a18_data_delayed_15 <= 0;
    a18_data_delayed_16 <= 0;
    a18_data_delayed_17 <= 0;
    a18_data_delayed_18 <= 0;
    a19_data_delayed_1 <= 0;
    a19_data_delayed_2 <= 0;
    a19_data_delayed_3 <= 0;
    a19_data_delayed_4 <= 0;
    a19_data_delayed_5 <= 0;
    a19_data_delayed_6 <= 0;
    a19_data_delayed_7 <= 0;
    a19_data_delayed_8 <= 0;
    a19_data_delayed_9 <= 0;
    a19_data_delayed_10 <= 0;
    a19_data_delayed_11 <= 0;
    a19_data_delayed_12 <= 0;
    a19_data_delayed_13 <= 0;
    a19_data_delayed_14 <= 0;
    a19_data_delayed_15 <= 0;
    a19_data_delayed_16 <= 0;
    a19_data_delayed_17 <= 0;
    a19_data_delayed_18 <= 0;
    a19_data_delayed_19 <= 0;
    a20_data_delayed_1 <= 0;
    a20_data_delayed_2 <= 0;
    a20_data_delayed_3 <= 0;
    a20_data_delayed_4 <= 0;
    a20_data_delayed_5 <= 0;
    a20_data_delayed_6 <= 0;
    a20_data_delayed_7 <= 0;
    a20_data_delayed_8 <= 0;
    a20_data_delayed_9 <= 0;
    a20_data_delayed_10 <= 0;
    a20_data_delayed_11 <= 0;
    a20_data_delayed_12 <= 0;
    a20_data_delayed_13 <= 0;
    a20_data_delayed_14 <= 0;
    a20_data_delayed_15 <= 0;
    a20_data_delayed_16 <= 0;
    a20_data_delayed_17 <= 0;
    a20_data_delayed_18 <= 0;
    a20_data_delayed_19 <= 0;
    a20_data_delayed_20 <= 0;
    a21_data_delayed_1 <= 0;
    a21_data_delayed_2 <= 0;
    a21_data_delayed_3 <= 0;
    a21_data_delayed_4 <= 0;
    a21_data_delayed_5 <= 0;
    a21_data_delayed_6 <= 0;
    a21_data_delayed_7 <= 0;
    a21_data_delayed_8 <= 0;
    a21_data_delayed_9 <= 0;
    a21_data_delayed_10 <= 0;
    a21_data_delayed_11 <= 0;
    a21_data_delayed_12 <= 0;
    a21_data_delayed_13 <= 0;
    a21_data_delayed_14 <= 0;
    a21_data_delayed_15 <= 0;
    a21_data_delayed_16 <= 0;
    a21_data_delayed_17 <= 0;
    a21_data_delayed_18 <= 0;
    a21_data_delayed_19 <= 0;
    a21_data_delayed_20 <= 0;
    a21_data_delayed_21 <= 0;
    a22_data_delayed_1 <= 0;
    a22_data_delayed_2 <= 0;
    a22_data_delayed_3 <= 0;
    a22_data_delayed_4 <= 0;
    a22_data_delayed_5 <= 0;
    a22_data_delayed_6 <= 0;
    a22_data_delayed_7 <= 0;
    a22_data_delayed_8 <= 0;
    a22_data_delayed_9 <= 0;
    a22_data_delayed_10 <= 0;
    a22_data_delayed_11 <= 0;
    a22_data_delayed_12 <= 0;
    a22_data_delayed_13 <= 0;
    a22_data_delayed_14 <= 0;
    a22_data_delayed_15 <= 0;
    a22_data_delayed_16 <= 0;
    a22_data_delayed_17 <= 0;
    a22_data_delayed_18 <= 0;
    a22_data_delayed_19 <= 0;
    a22_data_delayed_20 <= 0;
    a22_data_delayed_21 <= 0;
    a22_data_delayed_22 <= 0;
    a23_data_delayed_1 <= 0;
    a23_data_delayed_2 <= 0;
    a23_data_delayed_3 <= 0;
    a23_data_delayed_4 <= 0;
    a23_data_delayed_5 <= 0;
    a23_data_delayed_6 <= 0;
    a23_data_delayed_7 <= 0;
    a23_data_delayed_8 <= 0;
    a23_data_delayed_9 <= 0;
    a23_data_delayed_10 <= 0;
    a23_data_delayed_11 <= 0;
    a23_data_delayed_12 <= 0;
    a23_data_delayed_13 <= 0;
    a23_data_delayed_14 <= 0;
    a23_data_delayed_15 <= 0;
    a23_data_delayed_16 <= 0;
    a23_data_delayed_17 <= 0;
    a23_data_delayed_18 <= 0;
    a23_data_delayed_19 <= 0;
    a23_data_delayed_20 <= 0;
    a23_data_delayed_21 <= 0;
    a23_data_delayed_22 <= 0;
    a23_data_delayed_23 <= 0;
    a24_data_delayed_1 <= 0;
    a24_data_delayed_2 <= 0;
    a24_data_delayed_3 <= 0;
    a24_data_delayed_4 <= 0;
    a24_data_delayed_5 <= 0;
    a24_data_delayed_6 <= 0;
    a24_data_delayed_7 <= 0;
    a24_data_delayed_8 <= 0;
    a24_data_delayed_9 <= 0;
    a24_data_delayed_10 <= 0;
    a24_data_delayed_11 <= 0;
    a24_data_delayed_12 <= 0;
    a24_data_delayed_13 <= 0;
    a24_data_delayed_14 <= 0;
    a24_data_delayed_15 <= 0;
    a24_data_delayed_16 <= 0;
    a24_data_delayed_17 <= 0;
    a24_data_delayed_18 <= 0;
    a24_data_delayed_19 <= 0;
    a24_data_delayed_20 <= 0;
    a24_data_delayed_21 <= 0;
    a24_data_delayed_22 <= 0;
    a24_data_delayed_23 <= 0;
    a24_data_delayed_24 <= 0;
    a25_data_delayed_1 <= 0;
    a25_data_delayed_2 <= 0;
    a25_data_delayed_3 <= 0;
    a25_data_delayed_4 <= 0;
    a25_data_delayed_5 <= 0;
    a25_data_delayed_6 <= 0;
    a25_data_delayed_7 <= 0;
    a25_data_delayed_8 <= 0;
    a25_data_delayed_9 <= 0;
    a25_data_delayed_10 <= 0;
    a25_data_delayed_11 <= 0;
    a25_data_delayed_12 <= 0;
    a25_data_delayed_13 <= 0;
    a25_data_delayed_14 <= 0;
    a25_data_delayed_15 <= 0;
    a25_data_delayed_16 <= 0;
    a25_data_delayed_17 <= 0;
    a25_data_delayed_18 <= 0;
    a25_data_delayed_19 <= 0;
    a25_data_delayed_20 <= 0;
    a25_data_delayed_21 <= 0;
    a25_data_delayed_22 <= 0;
    a25_data_delayed_23 <= 0;
    a25_data_delayed_24 <= 0;
    a25_data_delayed_25 <= 0;
    a26_data_delayed_1 <= 0;
    a26_data_delayed_2 <= 0;
    a26_data_delayed_3 <= 0;
    a26_data_delayed_4 <= 0;
    a26_data_delayed_5 <= 0;
    a26_data_delayed_6 <= 0;
    a26_data_delayed_7 <= 0;
    a26_data_delayed_8 <= 0;
    a26_data_delayed_9 <= 0;
    a26_data_delayed_10 <= 0;
    a26_data_delayed_11 <= 0;
    a26_data_delayed_12 <= 0;
    a26_data_delayed_13 <= 0;
    a26_data_delayed_14 <= 0;
    a26_data_delayed_15 <= 0;
    a26_data_delayed_16 <= 0;
    a26_data_delayed_17 <= 0;
    a26_data_delayed_18 <= 0;
    a26_data_delayed_19 <= 0;
    a26_data_delayed_20 <= 0;
    a26_data_delayed_21 <= 0;
    a26_data_delayed_22 <= 0;
    a26_data_delayed_23 <= 0;
    a26_data_delayed_24 <= 0;
    a26_data_delayed_25 <= 0;
    a26_data_delayed_26 <= 0;
    a27_data_delayed_1 <= 0;
    a27_data_delayed_2 <= 0;
    a27_data_delayed_3 <= 0;
    a27_data_delayed_4 <= 0;
    a27_data_delayed_5 <= 0;
    a27_data_delayed_6 <= 0;
    a27_data_delayed_7 <= 0;
    a27_data_delayed_8 <= 0;
    a27_data_delayed_9 <= 0;
    a27_data_delayed_10 <= 0;
    a27_data_delayed_11 <= 0;
    a27_data_delayed_12 <= 0;
    a27_data_delayed_13 <= 0;
    a27_data_delayed_14 <= 0;
    a27_data_delayed_15 <= 0;
    a27_data_delayed_16 <= 0;
    a27_data_delayed_17 <= 0;
    a27_data_delayed_18 <= 0;
    a27_data_delayed_19 <= 0;
    a27_data_delayed_20 <= 0;
    a27_data_delayed_21 <= 0;
    a27_data_delayed_22 <= 0;
    a27_data_delayed_23 <= 0;
    a27_data_delayed_24 <= 0;
    a27_data_delayed_25 <= 0;
    a27_data_delayed_26 <= 0;
    a27_data_delayed_27 <= 0;
    a28_data_delayed_1 <= 0;
    a28_data_delayed_2 <= 0;
    a28_data_delayed_3 <= 0;
    a28_data_delayed_4 <= 0;
    a28_data_delayed_5 <= 0;
    a28_data_delayed_6 <= 0;
    a28_data_delayed_7 <= 0;
    a28_data_delayed_8 <= 0;
    a28_data_delayed_9 <= 0;
    a28_data_delayed_10 <= 0;
    a28_data_delayed_11 <= 0;
    a28_data_delayed_12 <= 0;
    a28_data_delayed_13 <= 0;
    a28_data_delayed_14 <= 0;
    a28_data_delayed_15 <= 0;
    a28_data_delayed_16 <= 0;
    a28_data_delayed_17 <= 0;
    a28_data_delayed_18 <= 0;
    a28_data_delayed_19 <= 0;
    a28_data_delayed_20 <= 0;
    a28_data_delayed_21 <= 0;
    a28_data_delayed_22 <= 0;
    a28_data_delayed_23 <= 0;
    a28_data_delayed_24 <= 0;
    a28_data_delayed_25 <= 0;
    a28_data_delayed_26 <= 0;
    a28_data_delayed_27 <= 0;
    a28_data_delayed_28 <= 0;
    a29_data_delayed_1 <= 0;
    a29_data_delayed_2 <= 0;
    a29_data_delayed_3 <= 0;
    a29_data_delayed_4 <= 0;
    a29_data_delayed_5 <= 0;
    a29_data_delayed_6 <= 0;
    a29_data_delayed_7 <= 0;
    a29_data_delayed_8 <= 0;
    a29_data_delayed_9 <= 0;
    a29_data_delayed_10 <= 0;
    a29_data_delayed_11 <= 0;
    a29_data_delayed_12 <= 0;
    a29_data_delayed_13 <= 0;
    a29_data_delayed_14 <= 0;
    a29_data_delayed_15 <= 0;
    a29_data_delayed_16 <= 0;
    a29_data_delayed_17 <= 0;
    a29_data_delayed_18 <= 0;
    a29_data_delayed_19 <= 0;
    a29_data_delayed_20 <= 0;
    a29_data_delayed_21 <= 0;
    a29_data_delayed_22 <= 0;
    a29_data_delayed_23 <= 0;
    a29_data_delayed_24 <= 0;
    a29_data_delayed_25 <= 0;
    a29_data_delayed_26 <= 0;
    a29_data_delayed_27 <= 0;
    a29_data_delayed_28 <= 0;
    a29_data_delayed_29 <= 0;
    a30_data_delayed_1 <= 0;
    a30_data_delayed_2 <= 0;
    a30_data_delayed_3 <= 0;
    a30_data_delayed_4 <= 0;
    a30_data_delayed_5 <= 0;
    a30_data_delayed_6 <= 0;
    a30_data_delayed_7 <= 0;
    a30_data_delayed_8 <= 0;
    a30_data_delayed_9 <= 0;
    a30_data_delayed_10 <= 0;
    a30_data_delayed_11 <= 0;
    a30_data_delayed_12 <= 0;
    a30_data_delayed_13 <= 0;
    a30_data_delayed_14 <= 0;
    a30_data_delayed_15 <= 0;
    a30_data_delayed_16 <= 0;
    a30_data_delayed_17 <= 0;
    a30_data_delayed_18 <= 0;
    a30_data_delayed_19 <= 0;
    a30_data_delayed_20 <= 0;
    a30_data_delayed_21 <= 0;
    a30_data_delayed_22 <= 0;
    a30_data_delayed_23 <= 0;
    a30_data_delayed_24 <= 0;
    a30_data_delayed_25 <= 0;
    a30_data_delayed_26 <= 0;
    a30_data_delayed_27 <= 0;
    a30_data_delayed_28 <= 0;
    a30_data_delayed_29 <= 0;
    a30_data_delayed_30 <= 0;
    a31_data_delayed_1 <= 0;
    a31_data_delayed_2 <= 0;
    a31_data_delayed_3 <= 0;
    a31_data_delayed_4 <= 0;
    a31_data_delayed_5 <= 0;
    a31_data_delayed_6 <= 0;
    a31_data_delayed_7 <= 0;
    a31_data_delayed_8 <= 0;
    a31_data_delayed_9 <= 0;
    a31_data_delayed_10 <= 0;
    a31_data_delayed_11 <= 0;
    a31_data_delayed_12 <= 0;
    a31_data_delayed_13 <= 0;
    a31_data_delayed_14 <= 0;
    a31_data_delayed_15 <= 0;
    a31_data_delayed_16 <= 0;
    a31_data_delayed_17 <= 0;
    a31_data_delayed_18 <= 0;
    a31_data_delayed_19 <= 0;
    a31_data_delayed_20 <= 0;
    a31_data_delayed_21 <= 0;
    a31_data_delayed_22 <= 0;
    a31_data_delayed_23 <= 0;
    a31_data_delayed_24 <= 0;
    a31_data_delayed_25 <= 0;
    a31_data_delayed_26 <= 0;
    a31_data_delayed_27 <= 0;
    a31_data_delayed_28 <= 0;
    a31_data_delayed_29 <= 0;
    a31_data_delayed_30 <= 0;
    a31_data_delayed_31 <= 0;

  end
  else begin
  a1_data_delayed_1 <= a1_data;
  a2_data_delayed_1 <= a2_data;
  a3_data_delayed_1 <= a3_data;
  a4_data_delayed_1 <= a4_data;
  a5_data_delayed_1 <= a5_data;
  a6_data_delayed_1 <= a6_data;
  a7_data_delayed_1 <= a7_data;
  a8_data_delayed_1 <= a8_data;
  a9_data_delayed_1 <= a9_data;
  a10_data_delayed_1 <= a10_data;
  a11_data_delayed_1 <= a11_data;
  a12_data_delayed_1 <= a12_data;
  a13_data_delayed_1 <= a13_data;
  a14_data_delayed_1 <= a14_data;
  a15_data_delayed_1 <= a15_data;
  a16_data_delayed_1 <= a16_data;
  a17_data_delayed_1 <= a17_data;
  a18_data_delayed_1 <= a18_data;
  a19_data_delayed_1 <= a19_data;
  a20_data_delayed_1 <= a20_data;
  a21_data_delayed_1 <= a21_data;
  a22_data_delayed_1 <= a22_data;
  a23_data_delayed_1 <= a23_data;
  a24_data_delayed_1 <= a24_data;
  a25_data_delayed_1 <= a25_data;
  a26_data_delayed_1 <= a26_data;
  a27_data_delayed_1 <= a27_data;
  a28_data_delayed_1 <= a28_data;
  a29_data_delayed_1 <= a29_data;
  a30_data_delayed_1 <= a30_data;
  a31_data_delayed_1 <= a31_data;
  a2_data_delayed_2 <= a2_data_delayed_1;
  a3_data_delayed_2 <= a3_data_delayed_1;
  a3_data_delayed_3 <= a3_data_delayed_2;
  a4_data_delayed_2 <= a4_data_delayed_1;
  a4_data_delayed_3 <= a4_data_delayed_2;
  a4_data_delayed_4 <= a4_data_delayed_3;
  a5_data_delayed_2 <= a5_data_delayed_1;
  a5_data_delayed_3 <= a5_data_delayed_2;
  a5_data_delayed_4 <= a5_data_delayed_3;
  a5_data_delayed_5 <= a5_data_delayed_4;
  a6_data_delayed_2 <= a6_data_delayed_1;
  a6_data_delayed_3 <= a6_data_delayed_2;
  a6_data_delayed_4 <= a6_data_delayed_3;
  a6_data_delayed_5 <= a6_data_delayed_4;
  a6_data_delayed_6 <= a6_data_delayed_5;
  a7_data_delayed_2 <= a7_data_delayed_1;
  a7_data_delayed_3 <= a7_data_delayed_2;
  a7_data_delayed_4 <= a7_data_delayed_3;
  a7_data_delayed_5 <= a7_data_delayed_4;
  a7_data_delayed_6 <= a7_data_delayed_5;
  a7_data_delayed_7 <= a7_data_delayed_6;
  a8_data_delayed_2 <= a8_data_delayed_1;
  a8_data_delayed_3 <= a8_data_delayed_2;
  a8_data_delayed_4 <= a8_data_delayed_3;
  a8_data_delayed_5 <= a8_data_delayed_4;
  a8_data_delayed_6 <= a8_data_delayed_5;
  a8_data_delayed_7 <= a8_data_delayed_6;
  a8_data_delayed_8 <= a8_data_delayed_7;
  a9_data_delayed_2 <= a9_data_delayed_1;
  a9_data_delayed_3 <= a9_data_delayed_2;
  a9_data_delayed_4 <= a9_data_delayed_3;
  a9_data_delayed_5 <= a9_data_delayed_4;
  a9_data_delayed_6 <= a9_data_delayed_5;
  a9_data_delayed_7 <= a9_data_delayed_6;
  a9_data_delayed_8 <= a9_data_delayed_7;
  a9_data_delayed_9 <= a9_data_delayed_8;
  a10_data_delayed_2 <= a10_data_delayed_1;
  a10_data_delayed_3 <= a10_data_delayed_2;
  a10_data_delayed_4 <= a10_data_delayed_3;
  a10_data_delayed_5 <= a10_data_delayed_4;
  a10_data_delayed_6 <= a10_data_delayed_5;
  a10_data_delayed_7 <= a10_data_delayed_6;
  a10_data_delayed_8 <= a10_data_delayed_7;
  a10_data_delayed_9 <= a10_data_delayed_8;
  a10_data_delayed_10 <= a10_data_delayed_9;
  a11_data_delayed_2 <= a11_data_delayed_1;
  a11_data_delayed_3 <= a11_data_delayed_2;
  a11_data_delayed_4 <= a11_data_delayed_3;
  a11_data_delayed_5 <= a11_data_delayed_4;
  a11_data_delayed_6 <= a11_data_delayed_5;
  a11_data_delayed_7 <= a11_data_delayed_6;
  a11_data_delayed_8 <= a11_data_delayed_7;
  a11_data_delayed_9 <= a11_data_delayed_8;
  a11_data_delayed_10 <= a11_data_delayed_9;
  a11_data_delayed_11 <= a11_data_delayed_10;
  a12_data_delayed_2 <= a12_data_delayed_1;
  a12_data_delayed_3 <= a12_data_delayed_2;
  a12_data_delayed_4 <= a12_data_delayed_3;
  a12_data_delayed_5 <= a12_data_delayed_4;
  a12_data_delayed_6 <= a12_data_delayed_5;
  a12_data_delayed_7 <= a12_data_delayed_6;
  a12_data_delayed_8 <= a12_data_delayed_7;
  a12_data_delayed_9 <= a12_data_delayed_8;
  a12_data_delayed_10 <= a12_data_delayed_9;
  a12_data_delayed_11 <= a12_data_delayed_10;
  a12_data_delayed_12 <= a12_data_delayed_11;
  a13_data_delayed_2 <= a13_data_delayed_1;
  a13_data_delayed_3 <= a13_data_delayed_2;
  a13_data_delayed_4 <= a13_data_delayed_3;
  a13_data_delayed_5 <= a13_data_delayed_4;
  a13_data_delayed_6 <= a13_data_delayed_5;
  a13_data_delayed_7 <= a13_data_delayed_6;
  a13_data_delayed_8 <= a13_data_delayed_7;
  a13_data_delayed_9 <= a13_data_delayed_8;
  a13_data_delayed_10 <= a13_data_delayed_9;
  a13_data_delayed_11 <= a13_data_delayed_10;
  a13_data_delayed_12 <= a13_data_delayed_11;
  a13_data_delayed_13 <= a13_data_delayed_12;
  a14_data_delayed_2 <= a14_data_delayed_1;
  a14_data_delayed_3 <= a14_data_delayed_2;
  a14_data_delayed_4 <= a14_data_delayed_3;
  a14_data_delayed_5 <= a14_data_delayed_4;
  a14_data_delayed_6 <= a14_data_delayed_5;
  a14_data_delayed_7 <= a14_data_delayed_6;
  a14_data_delayed_8 <= a14_data_delayed_7;
  a14_data_delayed_9 <= a14_data_delayed_8;
  a14_data_delayed_10 <= a14_data_delayed_9;
  a14_data_delayed_11 <= a14_data_delayed_10;
  a14_data_delayed_12 <= a14_data_delayed_11;
  a14_data_delayed_13 <= a14_data_delayed_12;
  a14_data_delayed_14 <= a14_data_delayed_13;
  a15_data_delayed_2 <= a15_data_delayed_1;
  a15_data_delayed_3 <= a15_data_delayed_2;
  a15_data_delayed_4 <= a15_data_delayed_3;
  a15_data_delayed_5 <= a15_data_delayed_4;
  a15_data_delayed_6 <= a15_data_delayed_5;
  a15_data_delayed_7 <= a15_data_delayed_6;
  a15_data_delayed_8 <= a15_data_delayed_7;
  a15_data_delayed_9 <= a15_data_delayed_8;
  a15_data_delayed_10 <= a15_data_delayed_9;
  a15_data_delayed_11 <= a15_data_delayed_10;
  a15_data_delayed_12 <= a15_data_delayed_11;
  a15_data_delayed_13 <= a15_data_delayed_12;
  a15_data_delayed_14 <= a15_data_delayed_13;
  a15_data_delayed_15 <= a15_data_delayed_14;
  a16_data_delayed_2 <= a16_data_delayed_1;
  a16_data_delayed_3 <= a16_data_delayed_2;
  a16_data_delayed_4 <= a16_data_delayed_3;
  a16_data_delayed_5 <= a16_data_delayed_4;
  a16_data_delayed_6 <= a16_data_delayed_5;
  a16_data_delayed_7 <= a16_data_delayed_6;
  a16_data_delayed_8 <= a16_data_delayed_7;
  a16_data_delayed_9 <= a16_data_delayed_8;
  a16_data_delayed_10 <= a16_data_delayed_9;
  a16_data_delayed_11 <= a16_data_delayed_10;
  a16_data_delayed_12 <= a16_data_delayed_11;
  a16_data_delayed_13 <= a16_data_delayed_12;
  a16_data_delayed_14 <= a16_data_delayed_13;
  a16_data_delayed_15 <= a16_data_delayed_14;
  a16_data_delayed_16 <= a16_data_delayed_15;
  a17_data_delayed_2 <= a17_data_delayed_1;
  a17_data_delayed_3 <= a17_data_delayed_2;
  a17_data_delayed_4 <= a17_data_delayed_3;
  a17_data_delayed_5 <= a17_data_delayed_4;
  a17_data_delayed_6 <= a17_data_delayed_5;
  a17_data_delayed_7 <= a17_data_delayed_6;
  a17_data_delayed_8 <= a17_data_delayed_7;
  a17_data_delayed_9 <= a17_data_delayed_8;
  a17_data_delayed_10 <= a17_data_delayed_9;
  a17_data_delayed_11 <= a17_data_delayed_10;
  a17_data_delayed_12 <= a17_data_delayed_11;
  a17_data_delayed_13 <= a17_data_delayed_12;
  a17_data_delayed_14 <= a17_data_delayed_13;
  a17_data_delayed_15 <= a17_data_delayed_14;
  a17_data_delayed_16 <= a17_data_delayed_15;
  a17_data_delayed_17 <= a17_data_delayed_16;
  a18_data_delayed_2 <= a18_data_delayed_1;
  a18_data_delayed_3 <= a18_data_delayed_2;
  a18_data_delayed_4 <= a18_data_delayed_3;
  a18_data_delayed_5 <= a18_data_delayed_4;
  a18_data_delayed_6 <= a18_data_delayed_5;
  a18_data_delayed_7 <= a18_data_delayed_6;
  a18_data_delayed_8 <= a18_data_delayed_7;
  a18_data_delayed_9 <= a18_data_delayed_8;
  a18_data_delayed_10 <= a18_data_delayed_9;
  a18_data_delayed_11 <= a18_data_delayed_10;
  a18_data_delayed_12 <= a18_data_delayed_11;
  a18_data_delayed_13 <= a18_data_delayed_12;
  a18_data_delayed_14 <= a18_data_delayed_13;
  a18_data_delayed_15 <= a18_data_delayed_14;
  a18_data_delayed_16 <= a18_data_delayed_15;
  a18_data_delayed_17 <= a18_data_delayed_16;
  a18_data_delayed_18 <= a18_data_delayed_17;
  a19_data_delayed_2 <= a19_data_delayed_1;
  a19_data_delayed_3 <= a19_data_delayed_2;
  a19_data_delayed_4 <= a19_data_delayed_3;
  a19_data_delayed_5 <= a19_data_delayed_4;
  a19_data_delayed_6 <= a19_data_delayed_5;
  a19_data_delayed_7 <= a19_data_delayed_6;
  a19_data_delayed_8 <= a19_data_delayed_7;
  a19_data_delayed_9 <= a19_data_delayed_8;
  a19_data_delayed_10 <= a19_data_delayed_9;
  a19_data_delayed_11 <= a19_data_delayed_10;
  a19_data_delayed_12 <= a19_data_delayed_11;
  a19_data_delayed_13 <= a19_data_delayed_12;
  a19_data_delayed_14 <= a19_data_delayed_13;
  a19_data_delayed_15 <= a19_data_delayed_14;
  a19_data_delayed_16 <= a19_data_delayed_15;
  a19_data_delayed_17 <= a19_data_delayed_16;
  a19_data_delayed_18 <= a19_data_delayed_17;
  a19_data_delayed_19 <= a19_data_delayed_18;
  a20_data_delayed_2 <= a20_data_delayed_1;
  a20_data_delayed_3 <= a20_data_delayed_2;
  a20_data_delayed_4 <= a20_data_delayed_3;
  a20_data_delayed_5 <= a20_data_delayed_4;
  a20_data_delayed_6 <= a20_data_delayed_5;
  a20_data_delayed_7 <= a20_data_delayed_6;
  a20_data_delayed_8 <= a20_data_delayed_7;
  a20_data_delayed_9 <= a20_data_delayed_8;
  a20_data_delayed_10 <= a20_data_delayed_9;
  a20_data_delayed_11 <= a20_data_delayed_10;
  a20_data_delayed_12 <= a20_data_delayed_11;
  a20_data_delayed_13 <= a20_data_delayed_12;
  a20_data_delayed_14 <= a20_data_delayed_13;
  a20_data_delayed_15 <= a20_data_delayed_14;
  a20_data_delayed_16 <= a20_data_delayed_15;
  a20_data_delayed_17 <= a20_data_delayed_16;
  a20_data_delayed_18 <= a20_data_delayed_17;
  a20_data_delayed_19 <= a20_data_delayed_18;
  a20_data_delayed_20 <= a20_data_delayed_19;
  a21_data_delayed_2 <= a21_data_delayed_1;
  a21_data_delayed_3 <= a21_data_delayed_2;
  a21_data_delayed_4 <= a21_data_delayed_3;
  a21_data_delayed_5 <= a21_data_delayed_4;
  a21_data_delayed_6 <= a21_data_delayed_5;
  a21_data_delayed_7 <= a21_data_delayed_6;
  a21_data_delayed_8 <= a21_data_delayed_7;
  a21_data_delayed_9 <= a21_data_delayed_8;
  a21_data_delayed_10 <= a21_data_delayed_9;
  a21_data_delayed_11 <= a21_data_delayed_10;
  a21_data_delayed_12 <= a21_data_delayed_11;
  a21_data_delayed_13 <= a21_data_delayed_12;
  a21_data_delayed_14 <= a21_data_delayed_13;
  a21_data_delayed_15 <= a21_data_delayed_14;
  a21_data_delayed_16 <= a21_data_delayed_15;
  a21_data_delayed_17 <= a21_data_delayed_16;
  a21_data_delayed_18 <= a21_data_delayed_17;
  a21_data_delayed_19 <= a21_data_delayed_18;
  a21_data_delayed_20 <= a21_data_delayed_19;
  a21_data_delayed_21 <= a21_data_delayed_20;
  a22_data_delayed_2 <= a22_data_delayed_1;
  a22_data_delayed_3 <= a22_data_delayed_2;
  a22_data_delayed_4 <= a22_data_delayed_3;
  a22_data_delayed_5 <= a22_data_delayed_4;
  a22_data_delayed_6 <= a22_data_delayed_5;
  a22_data_delayed_7 <= a22_data_delayed_6;
  a22_data_delayed_8 <= a22_data_delayed_7;
  a22_data_delayed_9 <= a22_data_delayed_8;
  a22_data_delayed_10 <= a22_data_delayed_9;
  a22_data_delayed_11 <= a22_data_delayed_10;
  a22_data_delayed_12 <= a22_data_delayed_11;
  a22_data_delayed_13 <= a22_data_delayed_12;
  a22_data_delayed_14 <= a22_data_delayed_13;
  a22_data_delayed_15 <= a22_data_delayed_14;
  a22_data_delayed_16 <= a22_data_delayed_15;
  a22_data_delayed_17 <= a22_data_delayed_16;
  a22_data_delayed_18 <= a22_data_delayed_17;
  a22_data_delayed_19 <= a22_data_delayed_18;
  a22_data_delayed_20 <= a22_data_delayed_19;
  a22_data_delayed_21 <= a22_data_delayed_20;
  a22_data_delayed_22 <= a22_data_delayed_21;
  a23_data_delayed_2 <= a23_data_delayed_1;
  a23_data_delayed_3 <= a23_data_delayed_2;
  a23_data_delayed_4 <= a23_data_delayed_3;
  a23_data_delayed_5 <= a23_data_delayed_4;
  a23_data_delayed_6 <= a23_data_delayed_5;
  a23_data_delayed_7 <= a23_data_delayed_6;
  a23_data_delayed_8 <= a23_data_delayed_7;
  a23_data_delayed_9 <= a23_data_delayed_8;
  a23_data_delayed_10 <= a23_data_delayed_9;
  a23_data_delayed_11 <= a23_data_delayed_10;
  a23_data_delayed_12 <= a23_data_delayed_11;
  a23_data_delayed_13 <= a23_data_delayed_12;
  a23_data_delayed_14 <= a23_data_delayed_13;
  a23_data_delayed_15 <= a23_data_delayed_14;
  a23_data_delayed_16 <= a23_data_delayed_15;
  a23_data_delayed_17 <= a23_data_delayed_16;
  a23_data_delayed_18 <= a23_data_delayed_17;
  a23_data_delayed_19 <= a23_data_delayed_18;
  a23_data_delayed_20 <= a23_data_delayed_19;
  a23_data_delayed_21 <= a23_data_delayed_20;
  a23_data_delayed_22 <= a23_data_delayed_21;
  a23_data_delayed_23 <= a23_data_delayed_22;
  a24_data_delayed_2 <= a24_data_delayed_1;
  a24_data_delayed_3 <= a24_data_delayed_2;
  a24_data_delayed_4 <= a24_data_delayed_3;
  a24_data_delayed_5 <= a24_data_delayed_4;
  a24_data_delayed_6 <= a24_data_delayed_5;
  a24_data_delayed_7 <= a24_data_delayed_6;
  a24_data_delayed_8 <= a24_data_delayed_7;
  a24_data_delayed_9 <= a24_data_delayed_8;
  a24_data_delayed_10 <= a24_data_delayed_9;
  a24_data_delayed_11 <= a24_data_delayed_10;
  a24_data_delayed_12 <= a24_data_delayed_11;
  a24_data_delayed_13 <= a24_data_delayed_12;
  a24_data_delayed_14 <= a24_data_delayed_13;
  a24_data_delayed_15 <= a24_data_delayed_14;
  a24_data_delayed_16 <= a24_data_delayed_15;
  a24_data_delayed_17 <= a24_data_delayed_16;
  a24_data_delayed_18 <= a24_data_delayed_17;
  a24_data_delayed_19 <= a24_data_delayed_18;
  a24_data_delayed_20 <= a24_data_delayed_19;
  a24_data_delayed_21 <= a24_data_delayed_20;
  a24_data_delayed_22 <= a24_data_delayed_21;
  a24_data_delayed_23 <= a24_data_delayed_22;
  a24_data_delayed_24 <= a24_data_delayed_23;
  a25_data_delayed_2 <= a25_data_delayed_1;
  a25_data_delayed_3 <= a25_data_delayed_2;
  a25_data_delayed_4 <= a25_data_delayed_3;
  a25_data_delayed_5 <= a25_data_delayed_4;
  a25_data_delayed_6 <= a25_data_delayed_5;
  a25_data_delayed_7 <= a25_data_delayed_6;
  a25_data_delayed_8 <= a25_data_delayed_7;
  a25_data_delayed_9 <= a25_data_delayed_8;
  a25_data_delayed_10 <= a25_data_delayed_9;
  a25_data_delayed_11 <= a25_data_delayed_10;
  a25_data_delayed_12 <= a25_data_delayed_11;
  a25_data_delayed_13 <= a25_data_delayed_12;
  a25_data_delayed_14 <= a25_data_delayed_13;
  a25_data_delayed_15 <= a25_data_delayed_14;
  a25_data_delayed_16 <= a25_data_delayed_15;
  a25_data_delayed_17 <= a25_data_delayed_16;
  a25_data_delayed_18 <= a25_data_delayed_17;
  a25_data_delayed_19 <= a25_data_delayed_18;
  a25_data_delayed_20 <= a25_data_delayed_19;
  a25_data_delayed_21 <= a25_data_delayed_20;
  a25_data_delayed_22 <= a25_data_delayed_21;
  a25_data_delayed_23 <= a25_data_delayed_22;
  a25_data_delayed_24 <= a25_data_delayed_23;
  a25_data_delayed_25 <= a25_data_delayed_24;
  a26_data_delayed_2 <= a26_data_delayed_1;
  a26_data_delayed_3 <= a26_data_delayed_2;
  a26_data_delayed_4 <= a26_data_delayed_3;
  a26_data_delayed_5 <= a26_data_delayed_4;
  a26_data_delayed_6 <= a26_data_delayed_5;
  a26_data_delayed_7 <= a26_data_delayed_6;
  a26_data_delayed_8 <= a26_data_delayed_7;
  a26_data_delayed_9 <= a26_data_delayed_8;
  a26_data_delayed_10 <= a26_data_delayed_9;
  a26_data_delayed_11 <= a26_data_delayed_10;
  a26_data_delayed_12 <= a26_data_delayed_11;
  a26_data_delayed_13 <= a26_data_delayed_12;
  a26_data_delayed_14 <= a26_data_delayed_13;
  a26_data_delayed_15 <= a26_data_delayed_14;
  a26_data_delayed_16 <= a26_data_delayed_15;
  a26_data_delayed_17 <= a26_data_delayed_16;
  a26_data_delayed_18 <= a26_data_delayed_17;
  a26_data_delayed_19 <= a26_data_delayed_18;
  a26_data_delayed_20 <= a26_data_delayed_19;
  a26_data_delayed_21 <= a26_data_delayed_20;
  a26_data_delayed_22 <= a26_data_delayed_21;
  a26_data_delayed_23 <= a26_data_delayed_22;
  a26_data_delayed_24 <= a26_data_delayed_23;
  a26_data_delayed_25 <= a26_data_delayed_24;
  a26_data_delayed_26 <= a26_data_delayed_25;
  a27_data_delayed_2 <= a27_data_delayed_1;
  a27_data_delayed_3 <= a27_data_delayed_2;
  a27_data_delayed_4 <= a27_data_delayed_3;
  a27_data_delayed_5 <= a27_data_delayed_4;
  a27_data_delayed_6 <= a27_data_delayed_5;
  a27_data_delayed_7 <= a27_data_delayed_6;
  a27_data_delayed_8 <= a27_data_delayed_7;
  a27_data_delayed_9 <= a27_data_delayed_8;
  a27_data_delayed_10 <= a27_data_delayed_9;
  a27_data_delayed_11 <= a27_data_delayed_10;
  a27_data_delayed_12 <= a27_data_delayed_11;
  a27_data_delayed_13 <= a27_data_delayed_12;
  a27_data_delayed_14 <= a27_data_delayed_13;
  a27_data_delayed_15 <= a27_data_delayed_14;
  a27_data_delayed_16 <= a27_data_delayed_15;
  a27_data_delayed_17 <= a27_data_delayed_16;
  a27_data_delayed_18 <= a27_data_delayed_17;
  a27_data_delayed_19 <= a27_data_delayed_18;
  a27_data_delayed_20 <= a27_data_delayed_19;
  a27_data_delayed_21 <= a27_data_delayed_20;
  a27_data_delayed_22 <= a27_data_delayed_21;
  a27_data_delayed_23 <= a27_data_delayed_22;
  a27_data_delayed_24 <= a27_data_delayed_23;
  a27_data_delayed_25 <= a27_data_delayed_24;
  a27_data_delayed_26 <= a27_data_delayed_25;
  a27_data_delayed_27 <= a27_data_delayed_26;
  a28_data_delayed_2 <= a28_data_delayed_1;
  a28_data_delayed_3 <= a28_data_delayed_2;
  a28_data_delayed_4 <= a28_data_delayed_3;
  a28_data_delayed_5 <= a28_data_delayed_4;
  a28_data_delayed_6 <= a28_data_delayed_5;
  a28_data_delayed_7 <= a28_data_delayed_6;
  a28_data_delayed_8 <= a28_data_delayed_7;
  a28_data_delayed_9 <= a28_data_delayed_8;
  a28_data_delayed_10 <= a28_data_delayed_9;
  a28_data_delayed_11 <= a28_data_delayed_10;
  a28_data_delayed_12 <= a28_data_delayed_11;
  a28_data_delayed_13 <= a28_data_delayed_12;
  a28_data_delayed_14 <= a28_data_delayed_13;
  a28_data_delayed_15 <= a28_data_delayed_14;
  a28_data_delayed_16 <= a28_data_delayed_15;
  a28_data_delayed_17 <= a28_data_delayed_16;
  a28_data_delayed_18 <= a28_data_delayed_17;
  a28_data_delayed_19 <= a28_data_delayed_18;
  a28_data_delayed_20 <= a28_data_delayed_19;
  a28_data_delayed_21 <= a28_data_delayed_20;
  a28_data_delayed_22 <= a28_data_delayed_21;
  a28_data_delayed_23 <= a28_data_delayed_22;
  a28_data_delayed_24 <= a28_data_delayed_23;
  a28_data_delayed_25 <= a28_data_delayed_24;
  a28_data_delayed_26 <= a28_data_delayed_25;
  a28_data_delayed_27 <= a28_data_delayed_26;
  a28_data_delayed_28 <= a28_data_delayed_27;
  a29_data_delayed_2 <= a29_data_delayed_1;
  a29_data_delayed_3 <= a29_data_delayed_2;
  a29_data_delayed_4 <= a29_data_delayed_3;
  a29_data_delayed_5 <= a29_data_delayed_4;
  a29_data_delayed_6 <= a29_data_delayed_5;
  a29_data_delayed_7 <= a29_data_delayed_6;
  a29_data_delayed_8 <= a29_data_delayed_7;
  a29_data_delayed_9 <= a29_data_delayed_8;
  a29_data_delayed_10 <= a29_data_delayed_9;
  a29_data_delayed_11 <= a29_data_delayed_10;
  a29_data_delayed_12 <= a29_data_delayed_11;
  a29_data_delayed_13 <= a29_data_delayed_12;
  a29_data_delayed_14 <= a29_data_delayed_13;
  a29_data_delayed_15 <= a29_data_delayed_14;
  a29_data_delayed_16 <= a29_data_delayed_15;
  a29_data_delayed_17 <= a29_data_delayed_16;
  a29_data_delayed_18 <= a29_data_delayed_17;
  a29_data_delayed_19 <= a29_data_delayed_18;
  a29_data_delayed_20 <= a29_data_delayed_19;
  a29_data_delayed_21 <= a29_data_delayed_20;
  a29_data_delayed_22 <= a29_data_delayed_21;
  a29_data_delayed_23 <= a29_data_delayed_22;
  a29_data_delayed_24 <= a29_data_delayed_23;
  a29_data_delayed_25 <= a29_data_delayed_24;
  a29_data_delayed_26 <= a29_data_delayed_25;
  a29_data_delayed_27 <= a29_data_delayed_26;
  a29_data_delayed_28 <= a29_data_delayed_27;
  a29_data_delayed_29 <= a29_data_delayed_28;
  a30_data_delayed_2 <= a30_data_delayed_1;
  a30_data_delayed_3 <= a30_data_delayed_2;
  a30_data_delayed_4 <= a30_data_delayed_3;
  a30_data_delayed_5 <= a30_data_delayed_4;
  a30_data_delayed_6 <= a30_data_delayed_5;
  a30_data_delayed_7 <= a30_data_delayed_6;
  a30_data_delayed_8 <= a30_data_delayed_7;
  a30_data_delayed_9 <= a30_data_delayed_8;
  a30_data_delayed_10 <= a30_data_delayed_9;
  a30_data_delayed_11 <= a30_data_delayed_10;
  a30_data_delayed_12 <= a30_data_delayed_11;
  a30_data_delayed_13 <= a30_data_delayed_12;
  a30_data_delayed_14 <= a30_data_delayed_13;
  a30_data_delayed_15 <= a30_data_delayed_14;
  a30_data_delayed_16 <= a30_data_delayed_15;
  a30_data_delayed_17 <= a30_data_delayed_16;
  a30_data_delayed_18 <= a30_data_delayed_17;
  a30_data_delayed_19 <= a30_data_delayed_18;
  a30_data_delayed_20 <= a30_data_delayed_19;
  a30_data_delayed_21 <= a30_data_delayed_20;
  a30_data_delayed_22 <= a30_data_delayed_21;
  a30_data_delayed_23 <= a30_data_delayed_22;
  a30_data_delayed_24 <= a30_data_delayed_23;
  a30_data_delayed_25 <= a30_data_delayed_24;
  a30_data_delayed_26 <= a30_data_delayed_25;
  a30_data_delayed_27 <= a30_data_delayed_26;
  a30_data_delayed_28 <= a30_data_delayed_27;
  a30_data_delayed_29 <= a30_data_delayed_28;
  a30_data_delayed_30 <= a30_data_delayed_29;
  a31_data_delayed_2 <= a31_data_delayed_1;
  a31_data_delayed_3 <= a31_data_delayed_2;
  a31_data_delayed_4 <= a31_data_delayed_3;
  a31_data_delayed_5 <= a31_data_delayed_4;
  a31_data_delayed_6 <= a31_data_delayed_5;
  a31_data_delayed_7 <= a31_data_delayed_6;
  a31_data_delayed_8 <= a31_data_delayed_7;
  a31_data_delayed_9 <= a31_data_delayed_8;
  a31_data_delayed_10 <= a31_data_delayed_9;
  a31_data_delayed_11 <= a31_data_delayed_10;
  a31_data_delayed_12 <= a31_data_delayed_11;
  a31_data_delayed_13 <= a31_data_delayed_12;
  a31_data_delayed_14 <= a31_data_delayed_13;
  a31_data_delayed_15 <= a31_data_delayed_14;
  a31_data_delayed_16 <= a31_data_delayed_15;
  a31_data_delayed_17 <= a31_data_delayed_16;
  a31_data_delayed_18 <= a31_data_delayed_17;
  a31_data_delayed_19 <= a31_data_delayed_18;
  a31_data_delayed_20 <= a31_data_delayed_19;
  a31_data_delayed_21 <= a31_data_delayed_20;
  a31_data_delayed_22 <= a31_data_delayed_21;
  a31_data_delayed_23 <= a31_data_delayed_22;
  a31_data_delayed_24 <= a31_data_delayed_23;
  a31_data_delayed_25 <= a31_data_delayed_24;
  a31_data_delayed_26 <= a31_data_delayed_25;
  a31_data_delayed_27 <= a31_data_delayed_26;
  a31_data_delayed_28 <= a31_data_delayed_27;
  a31_data_delayed_29 <= a31_data_delayed_28;
  a31_data_delayed_30 <= a31_data_delayed_29;
  a31_data_delayed_31 <= a31_data_delayed_30;
 
  end
end

//////////////////////////////////////////////////////////////////////////
// Logic to generate addresses to BRAM B
//////////////////////////////////////////////////////////////////////////
reg [`AWIDTH-1:0] b_addr;
reg b_mem_access; //flag that tells whether the matmul is trying to access memory or not
always @(posedge clk) begin
  //else if (clk_cnt >= b_loc*`MAT_MUL_SIZE+final_mat_mul_size) begin
  //Writing the line above to avoid multiplication:

  if ((reset || ~start_mat_mul) || (clk_cnt >= (b_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin

      b_addr <= address_mat_b - address_stride_b;
  
    b_mem_access <= 0;
  end
  //else if ((clk_cnt >= b_loc*`MAT_MUL_SIZE) && (clk_cnt < b_loc*`MAT_MUL_SIZE+final_mat_mul_size)) begin
  //Writing the line above to avoid multiplication:

  else if ((clk_cnt >= (b_loc<<`LOG2_MAT_MUL_SIZE)) && (clk_cnt < (b_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin

      b_addr <= b_addr + address_stride_b;
  
    b_mem_access <= 1;
  end
end 

//////////////////////////////////////////////////////////////////////////
// Logic to generate valid signals for data coming from BRAM B
//////////////////////////////////////////////////////////////////////////
reg [7:0] b_mem_access_counter;
always @(posedge clk) begin
  if (reset || ~start_mat_mul) begin
    b_mem_access_counter <= 0;
  end
  else if (b_mem_access == 1) begin
    b_mem_access_counter <= b_mem_access_counter + 1;  
  end
  else begin
    b_mem_access_counter <= 0;
  end
end

wire b_data_valid; //flag that tells whether the data from memory is valid
assign b_data_valid = 
     ((validity_mask_a_cols_b_rows[0]==1'b0 && b_mem_access_counter==1) ||
      (validity_mask_a_cols_b_rows[1]==1'b0 && b_mem_access_counter==2) ||
      (validity_mask_a_cols_b_rows[2]==1'b0 && b_mem_access_counter==3) ||
      (validity_mask_a_cols_b_rows[3]==1'b0 && b_mem_access_counter==4) ||
      (validity_mask_a_cols_b_rows[4]==1'b0 && b_mem_access_counter==5) ||
      (validity_mask_a_cols_b_rows[5]==1'b0 && b_mem_access_counter==6) ||
      (validity_mask_a_cols_b_rows[6]==1'b0 && b_mem_access_counter==7) ||
      (validity_mask_a_cols_b_rows[7]==1'b0 && b_mem_access_counter==8) ||
      (validity_mask_a_cols_b_rows[8]==1'b0 && b_mem_access_counter==9) ||
      (validity_mask_a_cols_b_rows[9]==1'b0 && b_mem_access_counter==10) ||
      (validity_mask_a_cols_b_rows[10]==1'b0 && b_mem_access_counter==11) ||
      (validity_mask_a_cols_b_rows[11]==1'b0 && b_mem_access_counter==12) ||
      (validity_mask_a_cols_b_rows[12]==1'b0 && b_mem_access_counter==13) ||
      (validity_mask_a_cols_b_rows[13]==1'b0 && b_mem_access_counter==14) ||
      (validity_mask_a_cols_b_rows[14]==1'b0 && b_mem_access_counter==15) ||
      (validity_mask_a_cols_b_rows[15]==1'b0 && b_mem_access_counter==16) ||
      (validity_mask_a_cols_b_rows[16]==1'b0 && b_mem_access_counter==17) ||
      (validity_mask_a_cols_b_rows[17]==1'b0 && b_mem_access_counter==18) ||
      (validity_mask_a_cols_b_rows[18]==1'b0 && b_mem_access_counter==19) ||
      (validity_mask_a_cols_b_rows[19]==1'b0 && b_mem_access_counter==20) ||
      (validity_mask_a_cols_b_rows[20]==1'b0 && b_mem_access_counter==21) ||
      (validity_mask_a_cols_b_rows[21]==1'b0 && b_mem_access_counter==22) ||
      (validity_mask_a_cols_b_rows[22]==1'b0 && b_mem_access_counter==23) ||
      (validity_mask_a_cols_b_rows[23]==1'b0 && b_mem_access_counter==24) ||
      (validity_mask_a_cols_b_rows[24]==1'b0 && b_mem_access_counter==25) ||
      (validity_mask_a_cols_b_rows[25]==1'b0 && b_mem_access_counter==26) ||
      (validity_mask_a_cols_b_rows[26]==1'b0 && b_mem_access_counter==27) ||
      (validity_mask_a_cols_b_rows[27]==1'b0 && b_mem_access_counter==28) ||
      (validity_mask_a_cols_b_rows[28]==1'b0 && b_mem_access_counter==29) ||
      (validity_mask_a_cols_b_rows[29]==1'b0 && b_mem_access_counter==30) ||
      (validity_mask_a_cols_b_rows[30]==1'b0 && b_mem_access_counter==31) ||
      (validity_mask_a_cols_b_rows[31]==1'b0 && b_mem_access_counter==32)) ?
    
        1'b0 : (b_mem_access_counter >= `MEM_ACCESS_LATENCY);

//////////////////////////////////////////////////////////////////////////
// Logic to delay certain parts of the data received from BRAM B (systolic data setup)
//////////////////////////////////////////////////////////////////////////
assign b0_data = b_data[1*`DWIDTH-1:0*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[0]}};
assign b1_data = b_data[2*`DWIDTH-1:1*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[1]}};
assign b2_data = b_data[3*`DWIDTH-1:2*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[2]}};
assign b3_data = b_data[4*`DWIDTH-1:3*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[3]}};
assign b4_data = b_data[5*`DWIDTH-1:4*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[4]}};
assign b5_data = b_data[6*`DWIDTH-1:5*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[5]}};
assign b6_data = b_data[7*`DWIDTH-1:6*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[6]}};
assign b7_data = b_data[8*`DWIDTH-1:7*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[7]}};
assign b8_data = b_data[9*`DWIDTH-1:8*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[8]}};
assign b9_data = b_data[10*`DWIDTH-1:9*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[9]}};
assign b10_data = b_data[11*`DWIDTH-1:10*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[10]}};
assign b11_data = b_data[12*`DWIDTH-1:11*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[11]}};
assign b12_data = b_data[13*`DWIDTH-1:12*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[12]}};
assign b13_data = b_data[14*`DWIDTH-1:13*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[13]}};
assign b14_data = b_data[15*`DWIDTH-1:14*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[14]}};
assign b15_data = b_data[16*`DWIDTH-1:15*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[15]}};
assign b16_data = b_data[17*`DWIDTH-1:16*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[16]}};
assign b17_data = b_data[18*`DWIDTH-1:17*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[17]}};
assign b18_data = b_data[19*`DWIDTH-1:18*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[18]}};
assign b19_data = b_data[20*`DWIDTH-1:19*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[19]}};
assign b20_data = b_data[21*`DWIDTH-1:20*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[20]}};
assign b21_data = b_data[22*`DWIDTH-1:21*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[21]}};
assign b22_data = b_data[23*`DWIDTH-1:22*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[22]}};
assign b23_data = b_data[24*`DWIDTH-1:23*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[23]}};
assign b24_data = b_data[25*`DWIDTH-1:24*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[24]}};
assign b25_data = b_data[26*`DWIDTH-1:25*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[25]}};
assign b26_data = b_data[27*`DWIDTH-1:26*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[26]}};
assign b27_data = b_data[28*`DWIDTH-1:27*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[27]}};
assign b28_data = b_data[29*`DWIDTH-1:28*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[28]}};
assign b29_data = b_data[30*`DWIDTH-1:29*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[29]}};
assign b30_data = b_data[31*`DWIDTH-1:30*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[30]}};
assign b31_data = b_data[32*`DWIDTH-1:31*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[31]}};

reg [`DWIDTH-1:0] b1_data_delayed_1;
reg [`DWIDTH-1:0] b2_data_delayed_1;
reg [`DWIDTH-1:0] b2_data_delayed_2;
reg [`DWIDTH-1:0] b3_data_delayed_1;
reg [`DWIDTH-1:0] b3_data_delayed_2;
reg [`DWIDTH-1:0] b3_data_delayed_3;
reg [`DWIDTH-1:0] b4_data_delayed_1;
reg [`DWIDTH-1:0] b4_data_delayed_2;
reg [`DWIDTH-1:0] b4_data_delayed_3;
reg [`DWIDTH-1:0] b4_data_delayed_4;
reg [`DWIDTH-1:0] b5_data_delayed_1;
reg [`DWIDTH-1:0] b5_data_delayed_2;
reg [`DWIDTH-1:0] b5_data_delayed_3;
reg [`DWIDTH-1:0] b5_data_delayed_4;
reg [`DWIDTH-1:0] b5_data_delayed_5;
reg [`DWIDTH-1:0] b6_data_delayed_1;
reg [`DWIDTH-1:0] b6_data_delayed_2;
reg [`DWIDTH-1:0] b6_data_delayed_3;
reg [`DWIDTH-1:0] b6_data_delayed_4;
reg [`DWIDTH-1:0] b6_data_delayed_5;
reg [`DWIDTH-1:0] b6_data_delayed_6;
reg [`DWIDTH-1:0] b7_data_delayed_1;
reg [`DWIDTH-1:0] b7_data_delayed_2;
reg [`DWIDTH-1:0] b7_data_delayed_3;
reg [`DWIDTH-1:0] b7_data_delayed_4;
reg [`DWIDTH-1:0] b7_data_delayed_5;
reg [`DWIDTH-1:0] b7_data_delayed_6;
reg [`DWIDTH-1:0] b7_data_delayed_7;
reg [`DWIDTH-1:0] b8_data_delayed_1;
reg [`DWIDTH-1:0] b8_data_delayed_2;
reg [`DWIDTH-1:0] b8_data_delayed_3;
reg [`DWIDTH-1:0] b8_data_delayed_4;
reg [`DWIDTH-1:0] b8_data_delayed_5;
reg [`DWIDTH-1:0] b8_data_delayed_6;
reg [`DWIDTH-1:0] b8_data_delayed_7;
reg [`DWIDTH-1:0] b8_data_delayed_8;
reg [`DWIDTH-1:0] b9_data_delayed_1;
reg [`DWIDTH-1:0] b9_data_delayed_2;
reg [`DWIDTH-1:0] b9_data_delayed_3;
reg [`DWIDTH-1:0] b9_data_delayed_4;
reg [`DWIDTH-1:0] b9_data_delayed_5;
reg [`DWIDTH-1:0] b9_data_delayed_6;
reg [`DWIDTH-1:0] b9_data_delayed_7;
reg [`DWIDTH-1:0] b9_data_delayed_8;
reg [`DWIDTH-1:0] b9_data_delayed_9;
reg [`DWIDTH-1:0] b10_data_delayed_1;
reg [`DWIDTH-1:0] b10_data_delayed_2;
reg [`DWIDTH-1:0] b10_data_delayed_3;
reg [`DWIDTH-1:0] b10_data_delayed_4;
reg [`DWIDTH-1:0] b10_data_delayed_5;
reg [`DWIDTH-1:0] b10_data_delayed_6;
reg [`DWIDTH-1:0] b10_data_delayed_7;
reg [`DWIDTH-1:0] b10_data_delayed_8;
reg [`DWIDTH-1:0] b10_data_delayed_9;
reg [`DWIDTH-1:0] b10_data_delayed_10;
reg [`DWIDTH-1:0] b11_data_delayed_1;
reg [`DWIDTH-1:0] b11_data_delayed_2;
reg [`DWIDTH-1:0] b11_data_delayed_3;
reg [`DWIDTH-1:0] b11_data_delayed_4;
reg [`DWIDTH-1:0] b11_data_delayed_5;
reg [`DWIDTH-1:0] b11_data_delayed_6;
reg [`DWIDTH-1:0] b11_data_delayed_7;
reg [`DWIDTH-1:0] b11_data_delayed_8;
reg [`DWIDTH-1:0] b11_data_delayed_9;
reg [`DWIDTH-1:0] b11_data_delayed_10;
reg [`DWIDTH-1:0] b11_data_delayed_11;
reg [`DWIDTH-1:0] b12_data_delayed_1;
reg [`DWIDTH-1:0] b12_data_delayed_2;
reg [`DWIDTH-1:0] b12_data_delayed_3;
reg [`DWIDTH-1:0] b12_data_delayed_4;
reg [`DWIDTH-1:0] b12_data_delayed_5;
reg [`DWIDTH-1:0] b12_data_delayed_6;
reg [`DWIDTH-1:0] b12_data_delayed_7;
reg [`DWIDTH-1:0] b12_data_delayed_8;
reg [`DWIDTH-1:0] b12_data_delayed_9;
reg [`DWIDTH-1:0] b12_data_delayed_10;
reg [`DWIDTH-1:0] b12_data_delayed_11;
reg [`DWIDTH-1:0] b12_data_delayed_12;
reg [`DWIDTH-1:0] b13_data_delayed_1;
reg [`DWIDTH-1:0] b13_data_delayed_2;
reg [`DWIDTH-1:0] b13_data_delayed_3;
reg [`DWIDTH-1:0] b13_data_delayed_4;
reg [`DWIDTH-1:0] b13_data_delayed_5;
reg [`DWIDTH-1:0] b13_data_delayed_6;
reg [`DWIDTH-1:0] b13_data_delayed_7;
reg [`DWIDTH-1:0] b13_data_delayed_8;
reg [`DWIDTH-1:0] b13_data_delayed_9;
reg [`DWIDTH-1:0] b13_data_delayed_10;
reg [`DWIDTH-1:0] b13_data_delayed_11;
reg [`DWIDTH-1:0] b13_data_delayed_12;
reg [`DWIDTH-1:0] b13_data_delayed_13;
reg [`DWIDTH-1:0] b14_data_delayed_1;
reg [`DWIDTH-1:0] b14_data_delayed_2;
reg [`DWIDTH-1:0] b14_data_delayed_3;
reg [`DWIDTH-1:0] b14_data_delayed_4;
reg [`DWIDTH-1:0] b14_data_delayed_5;
reg [`DWIDTH-1:0] b14_data_delayed_6;
reg [`DWIDTH-1:0] b14_data_delayed_7;
reg [`DWIDTH-1:0] b14_data_delayed_8;
reg [`DWIDTH-1:0] b14_data_delayed_9;
reg [`DWIDTH-1:0] b14_data_delayed_10;
reg [`DWIDTH-1:0] b14_data_delayed_11;
reg [`DWIDTH-1:0] b14_data_delayed_12;
reg [`DWIDTH-1:0] b14_data_delayed_13;
reg [`DWIDTH-1:0] b14_data_delayed_14;
reg [`DWIDTH-1:0] b15_data_delayed_1;
reg [`DWIDTH-1:0] b15_data_delayed_2;
reg [`DWIDTH-1:0] b15_data_delayed_3;
reg [`DWIDTH-1:0] b15_data_delayed_4;
reg [`DWIDTH-1:0] b15_data_delayed_5;
reg [`DWIDTH-1:0] b15_data_delayed_6;
reg [`DWIDTH-1:0] b15_data_delayed_7;
reg [`DWIDTH-1:0] b15_data_delayed_8;
reg [`DWIDTH-1:0] b15_data_delayed_9;
reg [`DWIDTH-1:0] b15_data_delayed_10;
reg [`DWIDTH-1:0] b15_data_delayed_11;
reg [`DWIDTH-1:0] b15_data_delayed_12;
reg [`DWIDTH-1:0] b15_data_delayed_13;
reg [`DWIDTH-1:0] b15_data_delayed_14;
reg [`DWIDTH-1:0] b15_data_delayed_15;
reg [`DWIDTH-1:0] b16_data_delayed_1;
reg [`DWIDTH-1:0] b16_data_delayed_2;
reg [`DWIDTH-1:0] b16_data_delayed_3;
reg [`DWIDTH-1:0] b16_data_delayed_4;
reg [`DWIDTH-1:0] b16_data_delayed_5;
reg [`DWIDTH-1:0] b16_data_delayed_6;
reg [`DWIDTH-1:0] b16_data_delayed_7;
reg [`DWIDTH-1:0] b16_data_delayed_8;
reg [`DWIDTH-1:0] b16_data_delayed_9;
reg [`DWIDTH-1:0] b16_data_delayed_10;
reg [`DWIDTH-1:0] b16_data_delayed_11;
reg [`DWIDTH-1:0] b16_data_delayed_12;
reg [`DWIDTH-1:0] b16_data_delayed_13;
reg [`DWIDTH-1:0] b16_data_delayed_14;
reg [`DWIDTH-1:0] b16_data_delayed_15;
reg [`DWIDTH-1:0] b16_data_delayed_16;
reg [`DWIDTH-1:0] b17_data_delayed_1;
reg [`DWIDTH-1:0] b17_data_delayed_2;
reg [`DWIDTH-1:0] b17_data_delayed_3;
reg [`DWIDTH-1:0] b17_data_delayed_4;
reg [`DWIDTH-1:0] b17_data_delayed_5;
reg [`DWIDTH-1:0] b17_data_delayed_6;
reg [`DWIDTH-1:0] b17_data_delayed_7;
reg [`DWIDTH-1:0] b17_data_delayed_8;
reg [`DWIDTH-1:0] b17_data_delayed_9;
reg [`DWIDTH-1:0] b17_data_delayed_10;
reg [`DWIDTH-1:0] b17_data_delayed_11;
reg [`DWIDTH-1:0] b17_data_delayed_12;
reg [`DWIDTH-1:0] b17_data_delayed_13;
reg [`DWIDTH-1:0] b17_data_delayed_14;
reg [`DWIDTH-1:0] b17_data_delayed_15;
reg [`DWIDTH-1:0] b17_data_delayed_16;
reg [`DWIDTH-1:0] b17_data_delayed_17;
reg [`DWIDTH-1:0] b18_data_delayed_1;
reg [`DWIDTH-1:0] b18_data_delayed_2;
reg [`DWIDTH-1:0] b18_data_delayed_3;
reg [`DWIDTH-1:0] b18_data_delayed_4;
reg [`DWIDTH-1:0] b18_data_delayed_5;
reg [`DWIDTH-1:0] b18_data_delayed_6;
reg [`DWIDTH-1:0] b18_data_delayed_7;
reg [`DWIDTH-1:0] b18_data_delayed_8;
reg [`DWIDTH-1:0] b18_data_delayed_9;
reg [`DWIDTH-1:0] b18_data_delayed_10;
reg [`DWIDTH-1:0] b18_data_delayed_11;
reg [`DWIDTH-1:0] b18_data_delayed_12;
reg [`DWIDTH-1:0] b18_data_delayed_13;
reg [`DWIDTH-1:0] b18_data_delayed_14;
reg [`DWIDTH-1:0] b18_data_delayed_15;
reg [`DWIDTH-1:0] b18_data_delayed_16;
reg [`DWIDTH-1:0] b18_data_delayed_17;
reg [`DWIDTH-1:0] b18_data_delayed_18;
reg [`DWIDTH-1:0] b19_data_delayed_1;
reg [`DWIDTH-1:0] b19_data_delayed_2;
reg [`DWIDTH-1:0] b19_data_delayed_3;
reg [`DWIDTH-1:0] b19_data_delayed_4;
reg [`DWIDTH-1:0] b19_data_delayed_5;
reg [`DWIDTH-1:0] b19_data_delayed_6;
reg [`DWIDTH-1:0] b19_data_delayed_7;
reg [`DWIDTH-1:0] b19_data_delayed_8;
reg [`DWIDTH-1:0] b19_data_delayed_9;
reg [`DWIDTH-1:0] b19_data_delayed_10;
reg [`DWIDTH-1:0] b19_data_delayed_11;
reg [`DWIDTH-1:0] b19_data_delayed_12;
reg [`DWIDTH-1:0] b19_data_delayed_13;
reg [`DWIDTH-1:0] b19_data_delayed_14;
reg [`DWIDTH-1:0] b19_data_delayed_15;
reg [`DWIDTH-1:0] b19_data_delayed_16;
reg [`DWIDTH-1:0] b19_data_delayed_17;
reg [`DWIDTH-1:0] b19_data_delayed_18;
reg [`DWIDTH-1:0] b19_data_delayed_19;
reg [`DWIDTH-1:0] b20_data_delayed_1;
reg [`DWIDTH-1:0] b20_data_delayed_2;
reg [`DWIDTH-1:0] b20_data_delayed_3;
reg [`DWIDTH-1:0] b20_data_delayed_4;
reg [`DWIDTH-1:0] b20_data_delayed_5;
reg [`DWIDTH-1:0] b20_data_delayed_6;
reg [`DWIDTH-1:0] b20_data_delayed_7;
reg [`DWIDTH-1:0] b20_data_delayed_8;
reg [`DWIDTH-1:0] b20_data_delayed_9;
reg [`DWIDTH-1:0] b20_data_delayed_10;
reg [`DWIDTH-1:0] b20_data_delayed_11;
reg [`DWIDTH-1:0] b20_data_delayed_12;
reg [`DWIDTH-1:0] b20_data_delayed_13;
reg [`DWIDTH-1:0] b20_data_delayed_14;
reg [`DWIDTH-1:0] b20_data_delayed_15;
reg [`DWIDTH-1:0] b20_data_delayed_16;
reg [`DWIDTH-1:0] b20_data_delayed_17;
reg [`DWIDTH-1:0] b20_data_delayed_18;
reg [`DWIDTH-1:0] b20_data_delayed_19;
reg [`DWIDTH-1:0] b20_data_delayed_20;
reg [`DWIDTH-1:0] b21_data_delayed_1;
reg [`DWIDTH-1:0] b21_data_delayed_2;
reg [`DWIDTH-1:0] b21_data_delayed_3;
reg [`DWIDTH-1:0] b21_data_delayed_4;
reg [`DWIDTH-1:0] b21_data_delayed_5;
reg [`DWIDTH-1:0] b21_data_delayed_6;
reg [`DWIDTH-1:0] b21_data_delayed_7;
reg [`DWIDTH-1:0] b21_data_delayed_8;
reg [`DWIDTH-1:0] b21_data_delayed_9;
reg [`DWIDTH-1:0] b21_data_delayed_10;
reg [`DWIDTH-1:0] b21_data_delayed_11;
reg [`DWIDTH-1:0] b21_data_delayed_12;
reg [`DWIDTH-1:0] b21_data_delayed_13;
reg [`DWIDTH-1:0] b21_data_delayed_14;
reg [`DWIDTH-1:0] b21_data_delayed_15;
reg [`DWIDTH-1:0] b21_data_delayed_16;
reg [`DWIDTH-1:0] b21_data_delayed_17;
reg [`DWIDTH-1:0] b21_data_delayed_18;
reg [`DWIDTH-1:0] b21_data_delayed_19;
reg [`DWIDTH-1:0] b21_data_delayed_20;
reg [`DWIDTH-1:0] b21_data_delayed_21;
reg [`DWIDTH-1:0] b22_data_delayed_1;
reg [`DWIDTH-1:0] b22_data_delayed_2;
reg [`DWIDTH-1:0] b22_data_delayed_3;
reg [`DWIDTH-1:0] b22_data_delayed_4;
reg [`DWIDTH-1:0] b22_data_delayed_5;
reg [`DWIDTH-1:0] b22_data_delayed_6;
reg [`DWIDTH-1:0] b22_data_delayed_7;
reg [`DWIDTH-1:0] b22_data_delayed_8;
reg [`DWIDTH-1:0] b22_data_delayed_9;
reg [`DWIDTH-1:0] b22_data_delayed_10;
reg [`DWIDTH-1:0] b22_data_delayed_11;
reg [`DWIDTH-1:0] b22_data_delayed_12;
reg [`DWIDTH-1:0] b22_data_delayed_13;
reg [`DWIDTH-1:0] b22_data_delayed_14;
reg [`DWIDTH-1:0] b22_data_delayed_15;
reg [`DWIDTH-1:0] b22_data_delayed_16;
reg [`DWIDTH-1:0] b22_data_delayed_17;
reg [`DWIDTH-1:0] b22_data_delayed_18;
reg [`DWIDTH-1:0] b22_data_delayed_19;
reg [`DWIDTH-1:0] b22_data_delayed_20;
reg [`DWIDTH-1:0] b22_data_delayed_21;
reg [`DWIDTH-1:0] b22_data_delayed_22;
reg [`DWIDTH-1:0] b23_data_delayed_1;
reg [`DWIDTH-1:0] b23_data_delayed_2;
reg [`DWIDTH-1:0] b23_data_delayed_3;
reg [`DWIDTH-1:0] b23_data_delayed_4;
reg [`DWIDTH-1:0] b23_data_delayed_5;
reg [`DWIDTH-1:0] b23_data_delayed_6;
reg [`DWIDTH-1:0] b23_data_delayed_7;
reg [`DWIDTH-1:0] b23_data_delayed_8;
reg [`DWIDTH-1:0] b23_data_delayed_9;
reg [`DWIDTH-1:0] b23_data_delayed_10;
reg [`DWIDTH-1:0] b23_data_delayed_11;
reg [`DWIDTH-1:0] b23_data_delayed_12;
reg [`DWIDTH-1:0] b23_data_delayed_13;
reg [`DWIDTH-1:0] b23_data_delayed_14;
reg [`DWIDTH-1:0] b23_data_delayed_15;
reg [`DWIDTH-1:0] b23_data_delayed_16;
reg [`DWIDTH-1:0] b23_data_delayed_17;
reg [`DWIDTH-1:0] b23_data_delayed_18;
reg [`DWIDTH-1:0] b23_data_delayed_19;
reg [`DWIDTH-1:0] b23_data_delayed_20;
reg [`DWIDTH-1:0] b23_data_delayed_21;
reg [`DWIDTH-1:0] b23_data_delayed_22;
reg [`DWIDTH-1:0] b23_data_delayed_23;
reg [`DWIDTH-1:0] b24_data_delayed_1;
reg [`DWIDTH-1:0] b24_data_delayed_2;
reg [`DWIDTH-1:0] b24_data_delayed_3;
reg [`DWIDTH-1:0] b24_data_delayed_4;
reg [`DWIDTH-1:0] b24_data_delayed_5;
reg [`DWIDTH-1:0] b24_data_delayed_6;
reg [`DWIDTH-1:0] b24_data_delayed_7;
reg [`DWIDTH-1:0] b24_data_delayed_8;
reg [`DWIDTH-1:0] b24_data_delayed_9;
reg [`DWIDTH-1:0] b24_data_delayed_10;
reg [`DWIDTH-1:0] b24_data_delayed_11;
reg [`DWIDTH-1:0] b24_data_delayed_12;
reg [`DWIDTH-1:0] b24_data_delayed_13;
reg [`DWIDTH-1:0] b24_data_delayed_14;
reg [`DWIDTH-1:0] b24_data_delayed_15;
reg [`DWIDTH-1:0] b24_data_delayed_16;
reg [`DWIDTH-1:0] b24_data_delayed_17;
reg [`DWIDTH-1:0] b24_data_delayed_18;
reg [`DWIDTH-1:0] b24_data_delayed_19;
reg [`DWIDTH-1:0] b24_data_delayed_20;
reg [`DWIDTH-1:0] b24_data_delayed_21;
reg [`DWIDTH-1:0] b24_data_delayed_22;
reg [`DWIDTH-1:0] b24_data_delayed_23;
reg [`DWIDTH-1:0] b24_data_delayed_24;
reg [`DWIDTH-1:0] b25_data_delayed_1;
reg [`DWIDTH-1:0] b25_data_delayed_2;
reg [`DWIDTH-1:0] b25_data_delayed_3;
reg [`DWIDTH-1:0] b25_data_delayed_4;
reg [`DWIDTH-1:0] b25_data_delayed_5;
reg [`DWIDTH-1:0] b25_data_delayed_6;
reg [`DWIDTH-1:0] b25_data_delayed_7;
reg [`DWIDTH-1:0] b25_data_delayed_8;
reg [`DWIDTH-1:0] b25_data_delayed_9;
reg [`DWIDTH-1:0] b25_data_delayed_10;
reg [`DWIDTH-1:0] b25_data_delayed_11;
reg [`DWIDTH-1:0] b25_data_delayed_12;
reg [`DWIDTH-1:0] b25_data_delayed_13;
reg [`DWIDTH-1:0] b25_data_delayed_14;
reg [`DWIDTH-1:0] b25_data_delayed_15;
reg [`DWIDTH-1:0] b25_data_delayed_16;
reg [`DWIDTH-1:0] b25_data_delayed_17;
reg [`DWIDTH-1:0] b25_data_delayed_18;
reg [`DWIDTH-1:0] b25_data_delayed_19;
reg [`DWIDTH-1:0] b25_data_delayed_20;
reg [`DWIDTH-1:0] b25_data_delayed_21;
reg [`DWIDTH-1:0] b25_data_delayed_22;
reg [`DWIDTH-1:0] b25_data_delayed_23;
reg [`DWIDTH-1:0] b25_data_delayed_24;
reg [`DWIDTH-1:0] b25_data_delayed_25;
reg [`DWIDTH-1:0] b26_data_delayed_1;
reg [`DWIDTH-1:0] b26_data_delayed_2;
reg [`DWIDTH-1:0] b26_data_delayed_3;
reg [`DWIDTH-1:0] b26_data_delayed_4;
reg [`DWIDTH-1:0] b26_data_delayed_5;
reg [`DWIDTH-1:0] b26_data_delayed_6;
reg [`DWIDTH-1:0] b26_data_delayed_7;
reg [`DWIDTH-1:0] b26_data_delayed_8;
reg [`DWIDTH-1:0] b26_data_delayed_9;
reg [`DWIDTH-1:0] b26_data_delayed_10;
reg [`DWIDTH-1:0] b26_data_delayed_11;
reg [`DWIDTH-1:0] b26_data_delayed_12;
reg [`DWIDTH-1:0] b26_data_delayed_13;
reg [`DWIDTH-1:0] b26_data_delayed_14;
reg [`DWIDTH-1:0] b26_data_delayed_15;
reg [`DWIDTH-1:0] b26_data_delayed_16;
reg [`DWIDTH-1:0] b26_data_delayed_17;
reg [`DWIDTH-1:0] b26_data_delayed_18;
reg [`DWIDTH-1:0] b26_data_delayed_19;
reg [`DWIDTH-1:0] b26_data_delayed_20;
reg [`DWIDTH-1:0] b26_data_delayed_21;
reg [`DWIDTH-1:0] b26_data_delayed_22;
reg [`DWIDTH-1:0] b26_data_delayed_23;
reg [`DWIDTH-1:0] b26_data_delayed_24;
reg [`DWIDTH-1:0] b26_data_delayed_25;
reg [`DWIDTH-1:0] b26_data_delayed_26;
reg [`DWIDTH-1:0] b27_data_delayed_1;
reg [`DWIDTH-1:0] b27_data_delayed_2;
reg [`DWIDTH-1:0] b27_data_delayed_3;
reg [`DWIDTH-1:0] b27_data_delayed_4;
reg [`DWIDTH-1:0] b27_data_delayed_5;
reg [`DWIDTH-1:0] b27_data_delayed_6;
reg [`DWIDTH-1:0] b27_data_delayed_7;
reg [`DWIDTH-1:0] b27_data_delayed_8;
reg [`DWIDTH-1:0] b27_data_delayed_9;
reg [`DWIDTH-1:0] b27_data_delayed_10;
reg [`DWIDTH-1:0] b27_data_delayed_11;
reg [`DWIDTH-1:0] b27_data_delayed_12;
reg [`DWIDTH-1:0] b27_data_delayed_13;
reg [`DWIDTH-1:0] b27_data_delayed_14;
reg [`DWIDTH-1:0] b27_data_delayed_15;
reg [`DWIDTH-1:0] b27_data_delayed_16;
reg [`DWIDTH-1:0] b27_data_delayed_17;
reg [`DWIDTH-1:0] b27_data_delayed_18;
reg [`DWIDTH-1:0] b27_data_delayed_19;
reg [`DWIDTH-1:0] b27_data_delayed_20;
reg [`DWIDTH-1:0] b27_data_delayed_21;
reg [`DWIDTH-1:0] b27_data_delayed_22;
reg [`DWIDTH-1:0] b27_data_delayed_23;
reg [`DWIDTH-1:0] b27_data_delayed_24;
reg [`DWIDTH-1:0] b27_data_delayed_25;
reg [`DWIDTH-1:0] b27_data_delayed_26;
reg [`DWIDTH-1:0] b27_data_delayed_27;
reg [`DWIDTH-1:0] b28_data_delayed_1;
reg [`DWIDTH-1:0] b28_data_delayed_2;
reg [`DWIDTH-1:0] b28_data_delayed_3;
reg [`DWIDTH-1:0] b28_data_delayed_4;
reg [`DWIDTH-1:0] b28_data_delayed_5;
reg [`DWIDTH-1:0] b28_data_delayed_6;
reg [`DWIDTH-1:0] b28_data_delayed_7;
reg [`DWIDTH-1:0] b28_data_delayed_8;
reg [`DWIDTH-1:0] b28_data_delayed_9;
reg [`DWIDTH-1:0] b28_data_delayed_10;
reg [`DWIDTH-1:0] b28_data_delayed_11;
reg [`DWIDTH-1:0] b28_data_delayed_12;
reg [`DWIDTH-1:0] b28_data_delayed_13;
reg [`DWIDTH-1:0] b28_data_delayed_14;
reg [`DWIDTH-1:0] b28_data_delayed_15;
reg [`DWIDTH-1:0] b28_data_delayed_16;
reg [`DWIDTH-1:0] b28_data_delayed_17;
reg [`DWIDTH-1:0] b28_data_delayed_18;
reg [`DWIDTH-1:0] b28_data_delayed_19;
reg [`DWIDTH-1:0] b28_data_delayed_20;
reg [`DWIDTH-1:0] b28_data_delayed_21;
reg [`DWIDTH-1:0] b28_data_delayed_22;
reg [`DWIDTH-1:0] b28_data_delayed_23;
reg [`DWIDTH-1:0] b28_data_delayed_24;
reg [`DWIDTH-1:0] b28_data_delayed_25;
reg [`DWIDTH-1:0] b28_data_delayed_26;
reg [`DWIDTH-1:0] b28_data_delayed_27;
reg [`DWIDTH-1:0] b28_data_delayed_28;
reg [`DWIDTH-1:0] b29_data_delayed_1;
reg [`DWIDTH-1:0] b29_data_delayed_2;
reg [`DWIDTH-1:0] b29_data_delayed_3;
reg [`DWIDTH-1:0] b29_data_delayed_4;
reg [`DWIDTH-1:0] b29_data_delayed_5;
reg [`DWIDTH-1:0] b29_data_delayed_6;
reg [`DWIDTH-1:0] b29_data_delayed_7;
reg [`DWIDTH-1:0] b29_data_delayed_8;
reg [`DWIDTH-1:0] b29_data_delayed_9;
reg [`DWIDTH-1:0] b29_data_delayed_10;
reg [`DWIDTH-1:0] b29_data_delayed_11;
reg [`DWIDTH-1:0] b29_data_delayed_12;
reg [`DWIDTH-1:0] b29_data_delayed_13;
reg [`DWIDTH-1:0] b29_data_delayed_14;
reg [`DWIDTH-1:0] b29_data_delayed_15;
reg [`DWIDTH-1:0] b29_data_delayed_16;
reg [`DWIDTH-1:0] b29_data_delayed_17;
reg [`DWIDTH-1:0] b29_data_delayed_18;
reg [`DWIDTH-1:0] b29_data_delayed_19;
reg [`DWIDTH-1:0] b29_data_delayed_20;
reg [`DWIDTH-1:0] b29_data_delayed_21;
reg [`DWIDTH-1:0] b29_data_delayed_22;
reg [`DWIDTH-1:0] b29_data_delayed_23;
reg [`DWIDTH-1:0] b29_data_delayed_24;
reg [`DWIDTH-1:0] b29_data_delayed_25;
reg [`DWIDTH-1:0] b29_data_delayed_26;
reg [`DWIDTH-1:0] b29_data_delayed_27;
reg [`DWIDTH-1:0] b29_data_delayed_28;
reg [`DWIDTH-1:0] b29_data_delayed_29;
reg [`DWIDTH-1:0] b30_data_delayed_1;
reg [`DWIDTH-1:0] b30_data_delayed_2;
reg [`DWIDTH-1:0] b30_data_delayed_3;
reg [`DWIDTH-1:0] b30_data_delayed_4;
reg [`DWIDTH-1:0] b30_data_delayed_5;
reg [`DWIDTH-1:0] b30_data_delayed_6;
reg [`DWIDTH-1:0] b30_data_delayed_7;
reg [`DWIDTH-1:0] b30_data_delayed_8;
reg [`DWIDTH-1:0] b30_data_delayed_9;
reg [`DWIDTH-1:0] b30_data_delayed_10;
reg [`DWIDTH-1:0] b30_data_delayed_11;
reg [`DWIDTH-1:0] b30_data_delayed_12;
reg [`DWIDTH-1:0] b30_data_delayed_13;
reg [`DWIDTH-1:0] b30_data_delayed_14;
reg [`DWIDTH-1:0] b30_data_delayed_15;
reg [`DWIDTH-1:0] b30_data_delayed_16;
reg [`DWIDTH-1:0] b30_data_delayed_17;
reg [`DWIDTH-1:0] b30_data_delayed_18;
reg [`DWIDTH-1:0] b30_data_delayed_19;
reg [`DWIDTH-1:0] b30_data_delayed_20;
reg [`DWIDTH-1:0] b30_data_delayed_21;
reg [`DWIDTH-1:0] b30_data_delayed_22;
reg [`DWIDTH-1:0] b30_data_delayed_23;
reg [`DWIDTH-1:0] b30_data_delayed_24;
reg [`DWIDTH-1:0] b30_data_delayed_25;
reg [`DWIDTH-1:0] b30_data_delayed_26;
reg [`DWIDTH-1:0] b30_data_delayed_27;
reg [`DWIDTH-1:0] b30_data_delayed_28;
reg [`DWIDTH-1:0] b30_data_delayed_29;
reg [`DWIDTH-1:0] b30_data_delayed_30;
reg [`DWIDTH-1:0] b31_data_delayed_1;
reg [`DWIDTH-1:0] b31_data_delayed_2;
reg [`DWIDTH-1:0] b31_data_delayed_3;
reg [`DWIDTH-1:0] b31_data_delayed_4;
reg [`DWIDTH-1:0] b31_data_delayed_5;
reg [`DWIDTH-1:0] b31_data_delayed_6;
reg [`DWIDTH-1:0] b31_data_delayed_7;
reg [`DWIDTH-1:0] b31_data_delayed_8;
reg [`DWIDTH-1:0] b31_data_delayed_9;
reg [`DWIDTH-1:0] b31_data_delayed_10;
reg [`DWIDTH-1:0] b31_data_delayed_11;
reg [`DWIDTH-1:0] b31_data_delayed_12;
reg [`DWIDTH-1:0] b31_data_delayed_13;
reg [`DWIDTH-1:0] b31_data_delayed_14;
reg [`DWIDTH-1:0] b31_data_delayed_15;
reg [`DWIDTH-1:0] b31_data_delayed_16;
reg [`DWIDTH-1:0] b31_data_delayed_17;
reg [`DWIDTH-1:0] b31_data_delayed_18;
reg [`DWIDTH-1:0] b31_data_delayed_19;
reg [`DWIDTH-1:0] b31_data_delayed_20;
reg [`DWIDTH-1:0] b31_data_delayed_21;
reg [`DWIDTH-1:0] b31_data_delayed_22;
reg [`DWIDTH-1:0] b31_data_delayed_23;
reg [`DWIDTH-1:0] b31_data_delayed_24;
reg [`DWIDTH-1:0] b31_data_delayed_25;
reg [`DWIDTH-1:0] b31_data_delayed_26;
reg [`DWIDTH-1:0] b31_data_delayed_27;
reg [`DWIDTH-1:0] b31_data_delayed_28;
reg [`DWIDTH-1:0] b31_data_delayed_29;
reg [`DWIDTH-1:0] b31_data_delayed_30;
reg [`DWIDTH-1:0] b31_data_delayed_31;


always @(posedge clk) begin
  if (reset || ~start_mat_mul || clk_cnt==0) begin
    b1_data_delayed_1 <= 0;
    b2_data_delayed_1 <= 0;
    b2_data_delayed_2 <= 0;
    b3_data_delayed_1 <= 0;
    b3_data_delayed_2 <= 0;
    b3_data_delayed_3 <= 0;
    b4_data_delayed_1 <= 0;
    b4_data_delayed_2 <= 0;
    b4_data_delayed_3 <= 0;
    b4_data_delayed_4 <= 0;
    b5_data_delayed_1 <= 0;
    b5_data_delayed_2 <= 0;
    b5_data_delayed_3 <= 0;
    b5_data_delayed_4 <= 0;
    b5_data_delayed_5 <= 0;
    b6_data_delayed_1 <= 0;
    b6_data_delayed_2 <= 0;
    b6_data_delayed_3 <= 0;
    b6_data_delayed_4 <= 0;
    b6_data_delayed_5 <= 0;
    b6_data_delayed_6 <= 0;
    b7_data_delayed_1 <= 0;
    b7_data_delayed_2 <= 0;
    b7_data_delayed_3 <= 0;
    b7_data_delayed_4 <= 0;
    b7_data_delayed_5 <= 0;
    b7_data_delayed_6 <= 0;
    b7_data_delayed_7 <= 0;
    b8_data_delayed_1 <= 0;
    b8_data_delayed_2 <= 0;
    b8_data_delayed_3 <= 0;
    b8_data_delayed_4 <= 0;
    b8_data_delayed_5 <= 0;
    b8_data_delayed_6 <= 0;
    b8_data_delayed_7 <= 0;
    b8_data_delayed_8 <= 0;
    b9_data_delayed_1 <= 0;
    b9_data_delayed_2 <= 0;
    b9_data_delayed_3 <= 0;
    b9_data_delayed_4 <= 0;
    b9_data_delayed_5 <= 0;
    b9_data_delayed_6 <= 0;
    b9_data_delayed_7 <= 0;
    b9_data_delayed_8 <= 0;
    b9_data_delayed_9 <= 0;
    b10_data_delayed_1 <= 0;
    b10_data_delayed_2 <= 0;
    b10_data_delayed_3 <= 0;
    b10_data_delayed_4 <= 0;
    b10_data_delayed_5 <= 0;
    b10_data_delayed_6 <= 0;
    b10_data_delayed_7 <= 0;
    b10_data_delayed_8 <= 0;
    b10_data_delayed_9 <= 0;
    b10_data_delayed_10 <= 0;
    b11_data_delayed_1 <= 0;
    b11_data_delayed_2 <= 0;
    b11_data_delayed_3 <= 0;
    b11_data_delayed_4 <= 0;
    b11_data_delayed_5 <= 0;
    b11_data_delayed_6 <= 0;
    b11_data_delayed_7 <= 0;
    b11_data_delayed_8 <= 0;
    b11_data_delayed_9 <= 0;
    b11_data_delayed_10 <= 0;
    b11_data_delayed_11 <= 0;
    b12_data_delayed_1 <= 0;
    b12_data_delayed_2 <= 0;
    b12_data_delayed_3 <= 0;
    b12_data_delayed_4 <= 0;
    b12_data_delayed_5 <= 0;
    b12_data_delayed_6 <= 0;
    b12_data_delayed_7 <= 0;
    b12_data_delayed_8 <= 0;
    b12_data_delayed_9 <= 0;
    b12_data_delayed_10 <= 0;
    b12_data_delayed_11 <= 0;
    b12_data_delayed_12 <= 0;
    b13_data_delayed_1 <= 0;
    b13_data_delayed_2 <= 0;
    b13_data_delayed_3 <= 0;
    b13_data_delayed_4 <= 0;
    b13_data_delayed_5 <= 0;
    b13_data_delayed_6 <= 0;
    b13_data_delayed_7 <= 0;
    b13_data_delayed_8 <= 0;
    b13_data_delayed_9 <= 0;
    b13_data_delayed_10 <= 0;
    b13_data_delayed_11 <= 0;
    b13_data_delayed_12 <= 0;
    b13_data_delayed_13 <= 0;
    b14_data_delayed_1 <= 0;
    b14_data_delayed_2 <= 0;
    b14_data_delayed_3 <= 0;
    b14_data_delayed_4 <= 0;
    b14_data_delayed_5 <= 0;
    b14_data_delayed_6 <= 0;
    b14_data_delayed_7 <= 0;
    b14_data_delayed_8 <= 0;
    b14_data_delayed_9 <= 0;
    b14_data_delayed_10 <= 0;
    b14_data_delayed_11 <= 0;
    b14_data_delayed_12 <= 0;
    b14_data_delayed_13 <= 0;
    b14_data_delayed_14 <= 0;
    b15_data_delayed_1 <= 0;
    b15_data_delayed_2 <= 0;
    b15_data_delayed_3 <= 0;
    b15_data_delayed_4 <= 0;
    b15_data_delayed_5 <= 0;
    b15_data_delayed_6 <= 0;
    b15_data_delayed_7 <= 0;
    b15_data_delayed_8 <= 0;
    b15_data_delayed_9 <= 0;
    b15_data_delayed_10 <= 0;
    b15_data_delayed_11 <= 0;
    b15_data_delayed_12 <= 0;
    b15_data_delayed_13 <= 0;
    b15_data_delayed_14 <= 0;
    b15_data_delayed_15 <= 0;
    b16_data_delayed_1 <= 0;
    b16_data_delayed_2 <= 0;
    b16_data_delayed_3 <= 0;
    b16_data_delayed_4 <= 0;
    b16_data_delayed_5 <= 0;
    b16_data_delayed_6 <= 0;
    b16_data_delayed_7 <= 0;
    b16_data_delayed_8 <= 0;
    b16_data_delayed_9 <= 0;
    b16_data_delayed_10 <= 0;
    b16_data_delayed_11 <= 0;
    b16_data_delayed_12 <= 0;
    b16_data_delayed_13 <= 0;
    b16_data_delayed_14 <= 0;
    b16_data_delayed_15 <= 0;
    b16_data_delayed_16 <= 0;
    b17_data_delayed_1 <= 0;
    b17_data_delayed_2 <= 0;
    b17_data_delayed_3 <= 0;
    b17_data_delayed_4 <= 0;
    b17_data_delayed_5 <= 0;
    b17_data_delayed_6 <= 0;
    b17_data_delayed_7 <= 0;
    b17_data_delayed_8 <= 0;
    b17_data_delayed_9 <= 0;
    b17_data_delayed_10 <= 0;
    b17_data_delayed_11 <= 0;
    b17_data_delayed_12 <= 0;
    b17_data_delayed_13 <= 0;
    b17_data_delayed_14 <= 0;
    b17_data_delayed_15 <= 0;
    b17_data_delayed_16 <= 0;
    b17_data_delayed_17 <= 0;
    b18_data_delayed_1 <= 0;
    b18_data_delayed_2 <= 0;
    b18_data_delayed_3 <= 0;
    b18_data_delayed_4 <= 0;
    b18_data_delayed_5 <= 0;
    b18_data_delayed_6 <= 0;
    b18_data_delayed_7 <= 0;
    b18_data_delayed_8 <= 0;
    b18_data_delayed_9 <= 0;
    b18_data_delayed_10 <= 0;
    b18_data_delayed_11 <= 0;
    b18_data_delayed_12 <= 0;
    b18_data_delayed_13 <= 0;
    b18_data_delayed_14 <= 0;
    b18_data_delayed_15 <= 0;
    b18_data_delayed_16 <= 0;
    b18_data_delayed_17 <= 0;
    b18_data_delayed_18 <= 0;
    b19_data_delayed_1 <= 0;
    b19_data_delayed_2 <= 0;
    b19_data_delayed_3 <= 0;
    b19_data_delayed_4 <= 0;
    b19_data_delayed_5 <= 0;
    b19_data_delayed_6 <= 0;
    b19_data_delayed_7 <= 0;
    b19_data_delayed_8 <= 0;
    b19_data_delayed_9 <= 0;
    b19_data_delayed_10 <= 0;
    b19_data_delayed_11 <= 0;
    b19_data_delayed_12 <= 0;
    b19_data_delayed_13 <= 0;
    b19_data_delayed_14 <= 0;
    b19_data_delayed_15 <= 0;
    b19_data_delayed_16 <= 0;
    b19_data_delayed_17 <= 0;
    b19_data_delayed_18 <= 0;
    b19_data_delayed_19 <= 0;
    b20_data_delayed_1 <= 0;
    b20_data_delayed_2 <= 0;
    b20_data_delayed_3 <= 0;
    b20_data_delayed_4 <= 0;
    b20_data_delayed_5 <= 0;
    b20_data_delayed_6 <= 0;
    b20_data_delayed_7 <= 0;
    b20_data_delayed_8 <= 0;
    b20_data_delayed_9 <= 0;
    b20_data_delayed_10 <= 0;
    b20_data_delayed_11 <= 0;
    b20_data_delayed_12 <= 0;
    b20_data_delayed_13 <= 0;
    b20_data_delayed_14 <= 0;
    b20_data_delayed_15 <= 0;
    b20_data_delayed_16 <= 0;
    b20_data_delayed_17 <= 0;
    b20_data_delayed_18 <= 0;
    b20_data_delayed_19 <= 0;
    b20_data_delayed_20 <= 0;
    b21_data_delayed_1 <= 0;
    b21_data_delayed_2 <= 0;
    b21_data_delayed_3 <= 0;
    b21_data_delayed_4 <= 0;
    b21_data_delayed_5 <= 0;
    b21_data_delayed_6 <= 0;
    b21_data_delayed_7 <= 0;
    b21_data_delayed_8 <= 0;
    b21_data_delayed_9 <= 0;
    b21_data_delayed_10 <= 0;
    b21_data_delayed_11 <= 0;
    b21_data_delayed_12 <= 0;
    b21_data_delayed_13 <= 0;
    b21_data_delayed_14 <= 0;
    b21_data_delayed_15 <= 0;
    b21_data_delayed_16 <= 0;
    b21_data_delayed_17 <= 0;
    b21_data_delayed_18 <= 0;
    b21_data_delayed_19 <= 0;
    b21_data_delayed_20 <= 0;
    b21_data_delayed_21 <= 0;
    b22_data_delayed_1 <= 0;
    b22_data_delayed_2 <= 0;
    b22_data_delayed_3 <= 0;
    b22_data_delayed_4 <= 0;
    b22_data_delayed_5 <= 0;
    b22_data_delayed_6 <= 0;
    b22_data_delayed_7 <= 0;
    b22_data_delayed_8 <= 0;
    b22_data_delayed_9 <= 0;
    b22_data_delayed_10 <= 0;
    b22_data_delayed_11 <= 0;
    b22_data_delayed_12 <= 0;
    b22_data_delayed_13 <= 0;
    b22_data_delayed_14 <= 0;
    b22_data_delayed_15 <= 0;
    b22_data_delayed_16 <= 0;
    b22_data_delayed_17 <= 0;
    b22_data_delayed_18 <= 0;
    b22_data_delayed_19 <= 0;
    b22_data_delayed_20 <= 0;
    b22_data_delayed_21 <= 0;
    b22_data_delayed_22 <= 0;
    b23_data_delayed_1 <= 0;
    b23_data_delayed_2 <= 0;
    b23_data_delayed_3 <= 0;
    b23_data_delayed_4 <= 0;
    b23_data_delayed_5 <= 0;
    b23_data_delayed_6 <= 0;
    b23_data_delayed_7 <= 0;
    b23_data_delayed_8 <= 0;
    b23_data_delayed_9 <= 0;
    b23_data_delayed_10 <= 0;
    b23_data_delayed_11 <= 0;
    b23_data_delayed_12 <= 0;
    b23_data_delayed_13 <= 0;
    b23_data_delayed_14 <= 0;
    b23_data_delayed_15 <= 0;
    b23_data_delayed_16 <= 0;
    b23_data_delayed_17 <= 0;
    b23_data_delayed_18 <= 0;
    b23_data_delayed_19 <= 0;
    b23_data_delayed_20 <= 0;
    b23_data_delayed_21 <= 0;
    b23_data_delayed_22 <= 0;
    b23_data_delayed_23 <= 0;
    b24_data_delayed_1 <= 0;
    b24_data_delayed_2 <= 0;
    b24_data_delayed_3 <= 0;
    b24_data_delayed_4 <= 0;
    b24_data_delayed_5 <= 0;
    b24_data_delayed_6 <= 0;
    b24_data_delayed_7 <= 0;
    b24_data_delayed_8 <= 0;
    b24_data_delayed_9 <= 0;
    b24_data_delayed_10 <= 0;
    b24_data_delayed_11 <= 0;
    b24_data_delayed_12 <= 0;
    b24_data_delayed_13 <= 0;
    b24_data_delayed_14 <= 0;
    b24_data_delayed_15 <= 0;
    b24_data_delayed_16 <= 0;
    b24_data_delayed_17 <= 0;
    b24_data_delayed_18 <= 0;
    b24_data_delayed_19 <= 0;
    b24_data_delayed_20 <= 0;
    b24_data_delayed_21 <= 0;
    b24_data_delayed_22 <= 0;
    b24_data_delayed_23 <= 0;
    b24_data_delayed_24 <= 0;
    b25_data_delayed_1 <= 0;
    b25_data_delayed_2 <= 0;
    b25_data_delayed_3 <= 0;
    b25_data_delayed_4 <= 0;
    b25_data_delayed_5 <= 0;
    b25_data_delayed_6 <= 0;
    b25_data_delayed_7 <= 0;
    b25_data_delayed_8 <= 0;
    b25_data_delayed_9 <= 0;
    b25_data_delayed_10 <= 0;
    b25_data_delayed_11 <= 0;
    b25_data_delayed_12 <= 0;
    b25_data_delayed_13 <= 0;
    b25_data_delayed_14 <= 0;
    b25_data_delayed_15 <= 0;
    b25_data_delayed_16 <= 0;
    b25_data_delayed_17 <= 0;
    b25_data_delayed_18 <= 0;
    b25_data_delayed_19 <= 0;
    b25_data_delayed_20 <= 0;
    b25_data_delayed_21 <= 0;
    b25_data_delayed_22 <= 0;
    b25_data_delayed_23 <= 0;
    b25_data_delayed_24 <= 0;
    b25_data_delayed_25 <= 0;
    b26_data_delayed_1 <= 0;
    b26_data_delayed_2 <= 0;
    b26_data_delayed_3 <= 0;
    b26_data_delayed_4 <= 0;
    b26_data_delayed_5 <= 0;
    b26_data_delayed_6 <= 0;
    b26_data_delayed_7 <= 0;
    b26_data_delayed_8 <= 0;
    b26_data_delayed_9 <= 0;
    b26_data_delayed_10 <= 0;
    b26_data_delayed_11 <= 0;
    b26_data_delayed_12 <= 0;
    b26_data_delayed_13 <= 0;
    b26_data_delayed_14 <= 0;
    b26_data_delayed_15 <= 0;
    b26_data_delayed_16 <= 0;
    b26_data_delayed_17 <= 0;
    b26_data_delayed_18 <= 0;
    b26_data_delayed_19 <= 0;
    b26_data_delayed_20 <= 0;
    b26_data_delayed_21 <= 0;
    b26_data_delayed_22 <= 0;
    b26_data_delayed_23 <= 0;
    b26_data_delayed_24 <= 0;
    b26_data_delayed_25 <= 0;
    b26_data_delayed_26 <= 0;
    b27_data_delayed_1 <= 0;
    b27_data_delayed_2 <= 0;
    b27_data_delayed_3 <= 0;
    b27_data_delayed_4 <= 0;
    b27_data_delayed_5 <= 0;
    b27_data_delayed_6 <= 0;
    b27_data_delayed_7 <= 0;
    b27_data_delayed_8 <= 0;
    b27_data_delayed_9 <= 0;
    b27_data_delayed_10 <= 0;
    b27_data_delayed_11 <= 0;
    b27_data_delayed_12 <= 0;
    b27_data_delayed_13 <= 0;
    b27_data_delayed_14 <= 0;
    b27_data_delayed_15 <= 0;
    b27_data_delayed_16 <= 0;
    b27_data_delayed_17 <= 0;
    b27_data_delayed_18 <= 0;
    b27_data_delayed_19 <= 0;
    b27_data_delayed_20 <= 0;
    b27_data_delayed_21 <= 0;
    b27_data_delayed_22 <= 0;
    b27_data_delayed_23 <= 0;
    b27_data_delayed_24 <= 0;
    b27_data_delayed_25 <= 0;
    b27_data_delayed_26 <= 0;
    b27_data_delayed_27 <= 0;
    b28_data_delayed_1 <= 0;
    b28_data_delayed_2 <= 0;
    b28_data_delayed_3 <= 0;
    b28_data_delayed_4 <= 0;
    b28_data_delayed_5 <= 0;
    b28_data_delayed_6 <= 0;
    b28_data_delayed_7 <= 0;
    b28_data_delayed_8 <= 0;
    b28_data_delayed_9 <= 0;
    b28_data_delayed_10 <= 0;
    b28_data_delayed_11 <= 0;
    b28_data_delayed_12 <= 0;
    b28_data_delayed_13 <= 0;
    b28_data_delayed_14 <= 0;
    b28_data_delayed_15 <= 0;
    b28_data_delayed_16 <= 0;
    b28_data_delayed_17 <= 0;
    b28_data_delayed_18 <= 0;
    b28_data_delayed_19 <= 0;
    b28_data_delayed_20 <= 0;
    b28_data_delayed_21 <= 0;
    b28_data_delayed_22 <= 0;
    b28_data_delayed_23 <= 0;
    b28_data_delayed_24 <= 0;
    b28_data_delayed_25 <= 0;
    b28_data_delayed_26 <= 0;
    b28_data_delayed_27 <= 0;
    b28_data_delayed_28 <= 0;
    b29_data_delayed_1 <= 0;
    b29_data_delayed_2 <= 0;
    b29_data_delayed_3 <= 0;
    b29_data_delayed_4 <= 0;
    b29_data_delayed_5 <= 0;
    b29_data_delayed_6 <= 0;
    b29_data_delayed_7 <= 0;
    b29_data_delayed_8 <= 0;
    b29_data_delayed_9 <= 0;
    b29_data_delayed_10 <= 0;
    b29_data_delayed_11 <= 0;
    b29_data_delayed_12 <= 0;
    b29_data_delayed_13 <= 0;
    b29_data_delayed_14 <= 0;
    b29_data_delayed_15 <= 0;
    b29_data_delayed_16 <= 0;
    b29_data_delayed_17 <= 0;
    b29_data_delayed_18 <= 0;
    b29_data_delayed_19 <= 0;
    b29_data_delayed_20 <= 0;
    b29_data_delayed_21 <= 0;
    b29_data_delayed_22 <= 0;
    b29_data_delayed_23 <= 0;
    b29_data_delayed_24 <= 0;
    b29_data_delayed_25 <= 0;
    b29_data_delayed_26 <= 0;
    b29_data_delayed_27 <= 0;
    b29_data_delayed_28 <= 0;
    b29_data_delayed_29 <= 0;
    b30_data_delayed_1 <= 0;
    b30_data_delayed_2 <= 0;
    b30_data_delayed_3 <= 0;
    b30_data_delayed_4 <= 0;
    b30_data_delayed_5 <= 0;
    b30_data_delayed_6 <= 0;
    b30_data_delayed_7 <= 0;
    b30_data_delayed_8 <= 0;
    b30_data_delayed_9 <= 0;
    b30_data_delayed_10 <= 0;
    b30_data_delayed_11 <= 0;
    b30_data_delayed_12 <= 0;
    b30_data_delayed_13 <= 0;
    b30_data_delayed_14 <= 0;
    b30_data_delayed_15 <= 0;
    b30_data_delayed_16 <= 0;
    b30_data_delayed_17 <= 0;
    b30_data_delayed_18 <= 0;
    b30_data_delayed_19 <= 0;
    b30_data_delayed_20 <= 0;
    b30_data_delayed_21 <= 0;
    b30_data_delayed_22 <= 0;
    b30_data_delayed_23 <= 0;
    b30_data_delayed_24 <= 0;
    b30_data_delayed_25 <= 0;
    b30_data_delayed_26 <= 0;
    b30_data_delayed_27 <= 0;
    b30_data_delayed_28 <= 0;
    b30_data_delayed_29 <= 0;
    b30_data_delayed_30 <= 0;
    b31_data_delayed_1 <= 0;
    b31_data_delayed_2 <= 0;
    b31_data_delayed_3 <= 0;
    b31_data_delayed_4 <= 0;
    b31_data_delayed_5 <= 0;
    b31_data_delayed_6 <= 0;
    b31_data_delayed_7 <= 0;
    b31_data_delayed_8 <= 0;
    b31_data_delayed_9 <= 0;
    b31_data_delayed_10 <= 0;
    b31_data_delayed_11 <= 0;
    b31_data_delayed_12 <= 0;
    b31_data_delayed_13 <= 0;
    b31_data_delayed_14 <= 0;
    b31_data_delayed_15 <= 0;
    b31_data_delayed_16 <= 0;
    b31_data_delayed_17 <= 0;
    b31_data_delayed_18 <= 0;
    b31_data_delayed_19 <= 0;
    b31_data_delayed_20 <= 0;
    b31_data_delayed_21 <= 0;
    b31_data_delayed_22 <= 0;
    b31_data_delayed_23 <= 0;
    b31_data_delayed_24 <= 0;
    b31_data_delayed_25 <= 0;
    b31_data_delayed_26 <= 0;
    b31_data_delayed_27 <= 0;
    b31_data_delayed_28 <= 0;
    b31_data_delayed_29 <= 0;
    b31_data_delayed_30 <= 0;
    b31_data_delayed_31 <= 0;

  end
  else begin
  b1_data_delayed_1 <= b1_data;
  b2_data_delayed_1 <= b2_data;
  b3_data_delayed_1 <= b3_data;
  b4_data_delayed_1 <= b4_data;
  b5_data_delayed_1 <= b5_data;
  b6_data_delayed_1 <= b6_data;
  b7_data_delayed_1 <= b7_data;
  b8_data_delayed_1 <= b8_data;
  b9_data_delayed_1 <= b9_data;
  b10_data_delayed_1 <= b10_data;
  b11_data_delayed_1 <= b11_data;
  b12_data_delayed_1 <= b12_data;
  b13_data_delayed_1 <= b13_data;
  b14_data_delayed_1 <= b14_data;
  b15_data_delayed_1 <= b15_data;
  b16_data_delayed_1 <= b16_data;
  b17_data_delayed_1 <= b17_data;
  b18_data_delayed_1 <= b18_data;
  b19_data_delayed_1 <= b19_data;
  b20_data_delayed_1 <= b20_data;
  b21_data_delayed_1 <= b21_data;
  b22_data_delayed_1 <= b22_data;
  b23_data_delayed_1 <= b23_data;
  b24_data_delayed_1 <= b24_data;
  b25_data_delayed_1 <= b25_data;
  b26_data_delayed_1 <= b26_data;
  b27_data_delayed_1 <= b27_data;
  b28_data_delayed_1 <= b28_data;
  b29_data_delayed_1 <= b29_data;
  b30_data_delayed_1 <= b30_data;
  b31_data_delayed_1 <= b31_data;
  b2_data_delayed_2 <= b2_data_delayed_1;
  b3_data_delayed_2 <= b3_data_delayed_1;
  b3_data_delayed_3 <= b3_data_delayed_2;
  b4_data_delayed_2 <= b4_data_delayed_1;
  b4_data_delayed_3 <= b4_data_delayed_2;
  b4_data_delayed_4 <= b4_data_delayed_3;
  b5_data_delayed_2 <= b5_data_delayed_1;
  b5_data_delayed_3 <= b5_data_delayed_2;
  b5_data_delayed_4 <= b5_data_delayed_3;
  b5_data_delayed_5 <= b5_data_delayed_4;
  b6_data_delayed_2 <= b6_data_delayed_1;
  b6_data_delayed_3 <= b6_data_delayed_2;
  b6_data_delayed_4 <= b6_data_delayed_3;
  b6_data_delayed_5 <= b6_data_delayed_4;
  b6_data_delayed_6 <= b6_data_delayed_5;
  b7_data_delayed_2 <= b7_data_delayed_1;
  b7_data_delayed_3 <= b7_data_delayed_2;
  b7_data_delayed_4 <= b7_data_delayed_3;
  b7_data_delayed_5 <= b7_data_delayed_4;
  b7_data_delayed_6 <= b7_data_delayed_5;
  b7_data_delayed_7 <= b7_data_delayed_6;
  b8_data_delayed_2 <= b8_data_delayed_1;
  b8_data_delayed_3 <= b8_data_delayed_2;
  b8_data_delayed_4 <= b8_data_delayed_3;
  b8_data_delayed_5 <= b8_data_delayed_4;
  b8_data_delayed_6 <= b8_data_delayed_5;
  b8_data_delayed_7 <= b8_data_delayed_6;
  b8_data_delayed_8 <= b8_data_delayed_7;
  b9_data_delayed_2 <= b9_data_delayed_1;
  b9_data_delayed_3 <= b9_data_delayed_2;
  b9_data_delayed_4 <= b9_data_delayed_3;
  b9_data_delayed_5 <= b9_data_delayed_4;
  b9_data_delayed_6 <= b9_data_delayed_5;
  b9_data_delayed_7 <= b9_data_delayed_6;
  b9_data_delayed_8 <= b9_data_delayed_7;
  b9_data_delayed_9 <= b9_data_delayed_8;
  b10_data_delayed_2 <= b10_data_delayed_1;
  b10_data_delayed_3 <= b10_data_delayed_2;
  b10_data_delayed_4 <= b10_data_delayed_3;
  b10_data_delayed_5 <= b10_data_delayed_4;
  b10_data_delayed_6 <= b10_data_delayed_5;
  b10_data_delayed_7 <= b10_data_delayed_6;
  b10_data_delayed_8 <= b10_data_delayed_7;
  b10_data_delayed_9 <= b10_data_delayed_8;
  b10_data_delayed_10 <= b10_data_delayed_9;
  b11_data_delayed_2 <= b11_data_delayed_1;
  b11_data_delayed_3 <= b11_data_delayed_2;
  b11_data_delayed_4 <= b11_data_delayed_3;
  b11_data_delayed_5 <= b11_data_delayed_4;
  b11_data_delayed_6 <= b11_data_delayed_5;
  b11_data_delayed_7 <= b11_data_delayed_6;
  b11_data_delayed_8 <= b11_data_delayed_7;
  b11_data_delayed_9 <= b11_data_delayed_8;
  b11_data_delayed_10 <= b11_data_delayed_9;
  b11_data_delayed_11 <= b11_data_delayed_10;
  b12_data_delayed_2 <= b12_data_delayed_1;
  b12_data_delayed_3 <= b12_data_delayed_2;
  b12_data_delayed_4 <= b12_data_delayed_3;
  b12_data_delayed_5 <= b12_data_delayed_4;
  b12_data_delayed_6 <= b12_data_delayed_5;
  b12_data_delayed_7 <= b12_data_delayed_6;
  b12_data_delayed_8 <= b12_data_delayed_7;
  b12_data_delayed_9 <= b12_data_delayed_8;
  b12_data_delayed_10 <= b12_data_delayed_9;
  b12_data_delayed_11 <= b12_data_delayed_10;
  b12_data_delayed_12 <= b12_data_delayed_11;
  b13_data_delayed_2 <= b13_data_delayed_1;
  b13_data_delayed_3 <= b13_data_delayed_2;
  b13_data_delayed_4 <= b13_data_delayed_3;
  b13_data_delayed_5 <= b13_data_delayed_4;
  b13_data_delayed_6 <= b13_data_delayed_5;
  b13_data_delayed_7 <= b13_data_delayed_6;
  b13_data_delayed_8 <= b13_data_delayed_7;
  b13_data_delayed_9 <= b13_data_delayed_8;
  b13_data_delayed_10 <= b13_data_delayed_9;
  b13_data_delayed_11 <= b13_data_delayed_10;
  b13_data_delayed_12 <= b13_data_delayed_11;
  b13_data_delayed_13 <= b13_data_delayed_12;
  b14_data_delayed_2 <= b14_data_delayed_1;
  b14_data_delayed_3 <= b14_data_delayed_2;
  b14_data_delayed_4 <= b14_data_delayed_3;
  b14_data_delayed_5 <= b14_data_delayed_4;
  b14_data_delayed_6 <= b14_data_delayed_5;
  b14_data_delayed_7 <= b14_data_delayed_6;
  b14_data_delayed_8 <= b14_data_delayed_7;
  b14_data_delayed_9 <= b14_data_delayed_8;
  b14_data_delayed_10 <= b14_data_delayed_9;
  b14_data_delayed_11 <= b14_data_delayed_10;
  b14_data_delayed_12 <= b14_data_delayed_11;
  b14_data_delayed_13 <= b14_data_delayed_12;
  b14_data_delayed_14 <= b14_data_delayed_13;
  b15_data_delayed_2 <= b15_data_delayed_1;
  b15_data_delayed_3 <= b15_data_delayed_2;
  b15_data_delayed_4 <= b15_data_delayed_3;
  b15_data_delayed_5 <= b15_data_delayed_4;
  b15_data_delayed_6 <= b15_data_delayed_5;
  b15_data_delayed_7 <= b15_data_delayed_6;
  b15_data_delayed_8 <= b15_data_delayed_7;
  b15_data_delayed_9 <= b15_data_delayed_8;
  b15_data_delayed_10 <= b15_data_delayed_9;
  b15_data_delayed_11 <= b15_data_delayed_10;
  b15_data_delayed_12 <= b15_data_delayed_11;
  b15_data_delayed_13 <= b15_data_delayed_12;
  b15_data_delayed_14 <= b15_data_delayed_13;
  b15_data_delayed_15 <= b15_data_delayed_14;
  b16_data_delayed_2 <= b16_data_delayed_1;
  b16_data_delayed_3 <= b16_data_delayed_2;
  b16_data_delayed_4 <= b16_data_delayed_3;
  b16_data_delayed_5 <= b16_data_delayed_4;
  b16_data_delayed_6 <= b16_data_delayed_5;
  b16_data_delayed_7 <= b16_data_delayed_6;
  b16_data_delayed_8 <= b16_data_delayed_7;
  b16_data_delayed_9 <= b16_data_delayed_8;
  b16_data_delayed_10 <= b16_data_delayed_9;
  b16_data_delayed_11 <= b16_data_delayed_10;
  b16_data_delayed_12 <= b16_data_delayed_11;
  b16_data_delayed_13 <= b16_data_delayed_12;
  b16_data_delayed_14 <= b16_data_delayed_13;
  b16_data_delayed_15 <= b16_data_delayed_14;
  b16_data_delayed_16 <= b16_data_delayed_15;
  b17_data_delayed_2 <= b17_data_delayed_1;
  b17_data_delayed_3 <= b17_data_delayed_2;
  b17_data_delayed_4 <= b17_data_delayed_3;
  b17_data_delayed_5 <= b17_data_delayed_4;
  b17_data_delayed_6 <= b17_data_delayed_5;
  b17_data_delayed_7 <= b17_data_delayed_6;
  b17_data_delayed_8 <= b17_data_delayed_7;
  b17_data_delayed_9 <= b17_data_delayed_8;
  b17_data_delayed_10 <= b17_data_delayed_9;
  b17_data_delayed_11 <= b17_data_delayed_10;
  b17_data_delayed_12 <= b17_data_delayed_11;
  b17_data_delayed_13 <= b17_data_delayed_12;
  b17_data_delayed_14 <= b17_data_delayed_13;
  b17_data_delayed_15 <= b17_data_delayed_14;
  b17_data_delayed_16 <= b17_data_delayed_15;
  b17_data_delayed_17 <= b17_data_delayed_16;
  b18_data_delayed_2 <= b18_data_delayed_1;
  b18_data_delayed_3 <= b18_data_delayed_2;
  b18_data_delayed_4 <= b18_data_delayed_3;
  b18_data_delayed_5 <= b18_data_delayed_4;
  b18_data_delayed_6 <= b18_data_delayed_5;
  b18_data_delayed_7 <= b18_data_delayed_6;
  b18_data_delayed_8 <= b18_data_delayed_7;
  b18_data_delayed_9 <= b18_data_delayed_8;
  b18_data_delayed_10 <= b18_data_delayed_9;
  b18_data_delayed_11 <= b18_data_delayed_10;
  b18_data_delayed_12 <= b18_data_delayed_11;
  b18_data_delayed_13 <= b18_data_delayed_12;
  b18_data_delayed_14 <= b18_data_delayed_13;
  b18_data_delayed_15 <= b18_data_delayed_14;
  b18_data_delayed_16 <= b18_data_delayed_15;
  b18_data_delayed_17 <= b18_data_delayed_16;
  b18_data_delayed_18 <= b18_data_delayed_17;
  b19_data_delayed_2 <= b19_data_delayed_1;
  b19_data_delayed_3 <= b19_data_delayed_2;
  b19_data_delayed_4 <= b19_data_delayed_3;
  b19_data_delayed_5 <= b19_data_delayed_4;
  b19_data_delayed_6 <= b19_data_delayed_5;
  b19_data_delayed_7 <= b19_data_delayed_6;
  b19_data_delayed_8 <= b19_data_delayed_7;
  b19_data_delayed_9 <= b19_data_delayed_8;
  b19_data_delayed_10 <= b19_data_delayed_9;
  b19_data_delayed_11 <= b19_data_delayed_10;
  b19_data_delayed_12 <= b19_data_delayed_11;
  b19_data_delayed_13 <= b19_data_delayed_12;
  b19_data_delayed_14 <= b19_data_delayed_13;
  b19_data_delayed_15 <= b19_data_delayed_14;
  b19_data_delayed_16 <= b19_data_delayed_15;
  b19_data_delayed_17 <= b19_data_delayed_16;
  b19_data_delayed_18 <= b19_data_delayed_17;
  b19_data_delayed_19 <= b19_data_delayed_18;
  b20_data_delayed_2 <= b20_data_delayed_1;
  b20_data_delayed_3 <= b20_data_delayed_2;
  b20_data_delayed_4 <= b20_data_delayed_3;
  b20_data_delayed_5 <= b20_data_delayed_4;
  b20_data_delayed_6 <= b20_data_delayed_5;
  b20_data_delayed_7 <= b20_data_delayed_6;
  b20_data_delayed_8 <= b20_data_delayed_7;
  b20_data_delayed_9 <= b20_data_delayed_8;
  b20_data_delayed_10 <= b20_data_delayed_9;
  b20_data_delayed_11 <= b20_data_delayed_10;
  b20_data_delayed_12 <= b20_data_delayed_11;
  b20_data_delayed_13 <= b20_data_delayed_12;
  b20_data_delayed_14 <= b20_data_delayed_13;
  b20_data_delayed_15 <= b20_data_delayed_14;
  b20_data_delayed_16 <= b20_data_delayed_15;
  b20_data_delayed_17 <= b20_data_delayed_16;
  b20_data_delayed_18 <= b20_data_delayed_17;
  b20_data_delayed_19 <= b20_data_delayed_18;
  b20_data_delayed_20 <= b20_data_delayed_19;
  b21_data_delayed_2 <= b21_data_delayed_1;
  b21_data_delayed_3 <= b21_data_delayed_2;
  b21_data_delayed_4 <= b21_data_delayed_3;
  b21_data_delayed_5 <= b21_data_delayed_4;
  b21_data_delayed_6 <= b21_data_delayed_5;
  b21_data_delayed_7 <= b21_data_delayed_6;
  b21_data_delayed_8 <= b21_data_delayed_7;
  b21_data_delayed_9 <= b21_data_delayed_8;
  b21_data_delayed_10 <= b21_data_delayed_9;
  b21_data_delayed_11 <= b21_data_delayed_10;
  b21_data_delayed_12 <= b21_data_delayed_11;
  b21_data_delayed_13 <= b21_data_delayed_12;
  b21_data_delayed_14 <= b21_data_delayed_13;
  b21_data_delayed_15 <= b21_data_delayed_14;
  b21_data_delayed_16 <= b21_data_delayed_15;
  b21_data_delayed_17 <= b21_data_delayed_16;
  b21_data_delayed_18 <= b21_data_delayed_17;
  b21_data_delayed_19 <= b21_data_delayed_18;
  b21_data_delayed_20 <= b21_data_delayed_19;
  b21_data_delayed_21 <= b21_data_delayed_20;
  b22_data_delayed_2 <= b22_data_delayed_1;
  b22_data_delayed_3 <= b22_data_delayed_2;
  b22_data_delayed_4 <= b22_data_delayed_3;
  b22_data_delayed_5 <= b22_data_delayed_4;
  b22_data_delayed_6 <= b22_data_delayed_5;
  b22_data_delayed_7 <= b22_data_delayed_6;
  b22_data_delayed_8 <= b22_data_delayed_7;
  b22_data_delayed_9 <= b22_data_delayed_8;
  b22_data_delayed_10 <= b22_data_delayed_9;
  b22_data_delayed_11 <= b22_data_delayed_10;
  b22_data_delayed_12 <= b22_data_delayed_11;
  b22_data_delayed_13 <= b22_data_delayed_12;
  b22_data_delayed_14 <= b22_data_delayed_13;
  b22_data_delayed_15 <= b22_data_delayed_14;
  b22_data_delayed_16 <= b22_data_delayed_15;
  b22_data_delayed_17 <= b22_data_delayed_16;
  b22_data_delayed_18 <= b22_data_delayed_17;
  b22_data_delayed_19 <= b22_data_delayed_18;
  b22_data_delayed_20 <= b22_data_delayed_19;
  b22_data_delayed_21 <= b22_data_delayed_20;
  b22_data_delayed_22 <= b22_data_delayed_21;
  b23_data_delayed_2 <= b23_data_delayed_1;
  b23_data_delayed_3 <= b23_data_delayed_2;
  b23_data_delayed_4 <= b23_data_delayed_3;
  b23_data_delayed_5 <= b23_data_delayed_4;
  b23_data_delayed_6 <= b23_data_delayed_5;
  b23_data_delayed_7 <= b23_data_delayed_6;
  b23_data_delayed_8 <= b23_data_delayed_7;
  b23_data_delayed_9 <= b23_data_delayed_8;
  b23_data_delayed_10 <= b23_data_delayed_9;
  b23_data_delayed_11 <= b23_data_delayed_10;
  b23_data_delayed_12 <= b23_data_delayed_11;
  b23_data_delayed_13 <= b23_data_delayed_12;
  b23_data_delayed_14 <= b23_data_delayed_13;
  b23_data_delayed_15 <= b23_data_delayed_14;
  b23_data_delayed_16 <= b23_data_delayed_15;
  b23_data_delayed_17 <= b23_data_delayed_16;
  b23_data_delayed_18 <= b23_data_delayed_17;
  b23_data_delayed_19 <= b23_data_delayed_18;
  b23_data_delayed_20 <= b23_data_delayed_19;
  b23_data_delayed_21 <= b23_data_delayed_20;
  b23_data_delayed_22 <= b23_data_delayed_21;
  b23_data_delayed_23 <= b23_data_delayed_22;
  b24_data_delayed_2 <= b24_data_delayed_1;
  b24_data_delayed_3 <= b24_data_delayed_2;
  b24_data_delayed_4 <= b24_data_delayed_3;
  b24_data_delayed_5 <= b24_data_delayed_4;
  b24_data_delayed_6 <= b24_data_delayed_5;
  b24_data_delayed_7 <= b24_data_delayed_6;
  b24_data_delayed_8 <= b24_data_delayed_7;
  b24_data_delayed_9 <= b24_data_delayed_8;
  b24_data_delayed_10 <= b24_data_delayed_9;
  b24_data_delayed_11 <= b24_data_delayed_10;
  b24_data_delayed_12 <= b24_data_delayed_11;
  b24_data_delayed_13 <= b24_data_delayed_12;
  b24_data_delayed_14 <= b24_data_delayed_13;
  b24_data_delayed_15 <= b24_data_delayed_14;
  b24_data_delayed_16 <= b24_data_delayed_15;
  b24_data_delayed_17 <= b24_data_delayed_16;
  b24_data_delayed_18 <= b24_data_delayed_17;
  b24_data_delayed_19 <= b24_data_delayed_18;
  b24_data_delayed_20 <= b24_data_delayed_19;
  b24_data_delayed_21 <= b24_data_delayed_20;
  b24_data_delayed_22 <= b24_data_delayed_21;
  b24_data_delayed_23 <= b24_data_delayed_22;
  b24_data_delayed_24 <= b24_data_delayed_23;
  b25_data_delayed_2 <= b25_data_delayed_1;
  b25_data_delayed_3 <= b25_data_delayed_2;
  b25_data_delayed_4 <= b25_data_delayed_3;
  b25_data_delayed_5 <= b25_data_delayed_4;
  b25_data_delayed_6 <= b25_data_delayed_5;
  b25_data_delayed_7 <= b25_data_delayed_6;
  b25_data_delayed_8 <= b25_data_delayed_7;
  b25_data_delayed_9 <= b25_data_delayed_8;
  b25_data_delayed_10 <= b25_data_delayed_9;
  b25_data_delayed_11 <= b25_data_delayed_10;
  b25_data_delayed_12 <= b25_data_delayed_11;
  b25_data_delayed_13 <= b25_data_delayed_12;
  b25_data_delayed_14 <= b25_data_delayed_13;
  b25_data_delayed_15 <= b25_data_delayed_14;
  b25_data_delayed_16 <= b25_data_delayed_15;
  b25_data_delayed_17 <= b25_data_delayed_16;
  b25_data_delayed_18 <= b25_data_delayed_17;
  b25_data_delayed_19 <= b25_data_delayed_18;
  b25_data_delayed_20 <= b25_data_delayed_19;
  b25_data_delayed_21 <= b25_data_delayed_20;
  b25_data_delayed_22 <= b25_data_delayed_21;
  b25_data_delayed_23 <= b25_data_delayed_22;
  b25_data_delayed_24 <= b25_data_delayed_23;
  b25_data_delayed_25 <= b25_data_delayed_24;
  b26_data_delayed_2 <= b26_data_delayed_1;
  b26_data_delayed_3 <= b26_data_delayed_2;
  b26_data_delayed_4 <= b26_data_delayed_3;
  b26_data_delayed_5 <= b26_data_delayed_4;
  b26_data_delayed_6 <= b26_data_delayed_5;
  b26_data_delayed_7 <= b26_data_delayed_6;
  b26_data_delayed_8 <= b26_data_delayed_7;
  b26_data_delayed_9 <= b26_data_delayed_8;
  b26_data_delayed_10 <= b26_data_delayed_9;
  b26_data_delayed_11 <= b26_data_delayed_10;
  b26_data_delayed_12 <= b26_data_delayed_11;
  b26_data_delayed_13 <= b26_data_delayed_12;
  b26_data_delayed_14 <= b26_data_delayed_13;
  b26_data_delayed_15 <= b26_data_delayed_14;
  b26_data_delayed_16 <= b26_data_delayed_15;
  b26_data_delayed_17 <= b26_data_delayed_16;
  b26_data_delayed_18 <= b26_data_delayed_17;
  b26_data_delayed_19 <= b26_data_delayed_18;
  b26_data_delayed_20 <= b26_data_delayed_19;
  b26_data_delayed_21 <= b26_data_delayed_20;
  b26_data_delayed_22 <= b26_data_delayed_21;
  b26_data_delayed_23 <= b26_data_delayed_22;
  b26_data_delayed_24 <= b26_data_delayed_23;
  b26_data_delayed_25 <= b26_data_delayed_24;
  b26_data_delayed_26 <= b26_data_delayed_25;
  b27_data_delayed_2 <= b27_data_delayed_1;
  b27_data_delayed_3 <= b27_data_delayed_2;
  b27_data_delayed_4 <= b27_data_delayed_3;
  b27_data_delayed_5 <= b27_data_delayed_4;
  b27_data_delayed_6 <= b27_data_delayed_5;
  b27_data_delayed_7 <= b27_data_delayed_6;
  b27_data_delayed_8 <= b27_data_delayed_7;
  b27_data_delayed_9 <= b27_data_delayed_8;
  b27_data_delayed_10 <= b27_data_delayed_9;
  b27_data_delayed_11 <= b27_data_delayed_10;
  b27_data_delayed_12 <= b27_data_delayed_11;
  b27_data_delayed_13 <= b27_data_delayed_12;
  b27_data_delayed_14 <= b27_data_delayed_13;
  b27_data_delayed_15 <= b27_data_delayed_14;
  b27_data_delayed_16 <= b27_data_delayed_15;
  b27_data_delayed_17 <= b27_data_delayed_16;
  b27_data_delayed_18 <= b27_data_delayed_17;
  b27_data_delayed_19 <= b27_data_delayed_18;
  b27_data_delayed_20 <= b27_data_delayed_19;
  b27_data_delayed_21 <= b27_data_delayed_20;
  b27_data_delayed_22 <= b27_data_delayed_21;
  b27_data_delayed_23 <= b27_data_delayed_22;
  b27_data_delayed_24 <= b27_data_delayed_23;
  b27_data_delayed_25 <= b27_data_delayed_24;
  b27_data_delayed_26 <= b27_data_delayed_25;
  b27_data_delayed_27 <= b27_data_delayed_26;
  b28_data_delayed_2 <= b28_data_delayed_1;
  b28_data_delayed_3 <= b28_data_delayed_2;
  b28_data_delayed_4 <= b28_data_delayed_3;
  b28_data_delayed_5 <= b28_data_delayed_4;
  b28_data_delayed_6 <= b28_data_delayed_5;
  b28_data_delayed_7 <= b28_data_delayed_6;
  b28_data_delayed_8 <= b28_data_delayed_7;
  b28_data_delayed_9 <= b28_data_delayed_8;
  b28_data_delayed_10 <= b28_data_delayed_9;
  b28_data_delayed_11 <= b28_data_delayed_10;
  b28_data_delayed_12 <= b28_data_delayed_11;
  b28_data_delayed_13 <= b28_data_delayed_12;
  b28_data_delayed_14 <= b28_data_delayed_13;
  b28_data_delayed_15 <= b28_data_delayed_14;
  b28_data_delayed_16 <= b28_data_delayed_15;
  b28_data_delayed_17 <= b28_data_delayed_16;
  b28_data_delayed_18 <= b28_data_delayed_17;
  b28_data_delayed_19 <= b28_data_delayed_18;
  b28_data_delayed_20 <= b28_data_delayed_19;
  b28_data_delayed_21 <= b28_data_delayed_20;
  b28_data_delayed_22 <= b28_data_delayed_21;
  b28_data_delayed_23 <= b28_data_delayed_22;
  b28_data_delayed_24 <= b28_data_delayed_23;
  b28_data_delayed_25 <= b28_data_delayed_24;
  b28_data_delayed_26 <= b28_data_delayed_25;
  b28_data_delayed_27 <= b28_data_delayed_26;
  b28_data_delayed_28 <= b28_data_delayed_27;
  b29_data_delayed_2 <= b29_data_delayed_1;
  b29_data_delayed_3 <= b29_data_delayed_2;
  b29_data_delayed_4 <= b29_data_delayed_3;
  b29_data_delayed_5 <= b29_data_delayed_4;
  b29_data_delayed_6 <= b29_data_delayed_5;
  b29_data_delayed_7 <= b29_data_delayed_6;
  b29_data_delayed_8 <= b29_data_delayed_7;
  b29_data_delayed_9 <= b29_data_delayed_8;
  b29_data_delayed_10 <= b29_data_delayed_9;
  b29_data_delayed_11 <= b29_data_delayed_10;
  b29_data_delayed_12 <= b29_data_delayed_11;
  b29_data_delayed_13 <= b29_data_delayed_12;
  b29_data_delayed_14 <= b29_data_delayed_13;
  b29_data_delayed_15 <= b29_data_delayed_14;
  b29_data_delayed_16 <= b29_data_delayed_15;
  b29_data_delayed_17 <= b29_data_delayed_16;
  b29_data_delayed_18 <= b29_data_delayed_17;
  b29_data_delayed_19 <= b29_data_delayed_18;
  b29_data_delayed_20 <= b29_data_delayed_19;
  b29_data_delayed_21 <= b29_data_delayed_20;
  b29_data_delayed_22 <= b29_data_delayed_21;
  b29_data_delayed_23 <= b29_data_delayed_22;
  b29_data_delayed_24 <= b29_data_delayed_23;
  b29_data_delayed_25 <= b29_data_delayed_24;
  b29_data_delayed_26 <= b29_data_delayed_25;
  b29_data_delayed_27 <= b29_data_delayed_26;
  b29_data_delayed_28 <= b29_data_delayed_27;
  b29_data_delayed_29 <= b29_data_delayed_28;
  b30_data_delayed_2 <= b30_data_delayed_1;
  b30_data_delayed_3 <= b30_data_delayed_2;
  b30_data_delayed_4 <= b30_data_delayed_3;
  b30_data_delayed_5 <= b30_data_delayed_4;
  b30_data_delayed_6 <= b30_data_delayed_5;
  b30_data_delayed_7 <= b30_data_delayed_6;
  b30_data_delayed_8 <= b30_data_delayed_7;
  b30_data_delayed_9 <= b30_data_delayed_8;
  b30_data_delayed_10 <= b30_data_delayed_9;
  b30_data_delayed_11 <= b30_data_delayed_10;
  b30_data_delayed_12 <= b30_data_delayed_11;
  b30_data_delayed_13 <= b30_data_delayed_12;
  b30_data_delayed_14 <= b30_data_delayed_13;
  b30_data_delayed_15 <= b30_data_delayed_14;
  b30_data_delayed_16 <= b30_data_delayed_15;
  b30_data_delayed_17 <= b30_data_delayed_16;
  b30_data_delayed_18 <= b30_data_delayed_17;
  b30_data_delayed_19 <= b30_data_delayed_18;
  b30_data_delayed_20 <= b30_data_delayed_19;
  b30_data_delayed_21 <= b30_data_delayed_20;
  b30_data_delayed_22 <= b30_data_delayed_21;
  b30_data_delayed_23 <= b30_data_delayed_22;
  b30_data_delayed_24 <= b30_data_delayed_23;
  b30_data_delayed_25 <= b30_data_delayed_24;
  b30_data_delayed_26 <= b30_data_delayed_25;
  b30_data_delayed_27 <= b30_data_delayed_26;
  b30_data_delayed_28 <= b30_data_delayed_27;
  b30_data_delayed_29 <= b30_data_delayed_28;
  b30_data_delayed_30 <= b30_data_delayed_29;
  b31_data_delayed_2 <= b31_data_delayed_1;
  b31_data_delayed_3 <= b31_data_delayed_2;
  b31_data_delayed_4 <= b31_data_delayed_3;
  b31_data_delayed_5 <= b31_data_delayed_4;
  b31_data_delayed_6 <= b31_data_delayed_5;
  b31_data_delayed_7 <= b31_data_delayed_6;
  b31_data_delayed_8 <= b31_data_delayed_7;
  b31_data_delayed_9 <= b31_data_delayed_8;
  b31_data_delayed_10 <= b31_data_delayed_9;
  b31_data_delayed_11 <= b31_data_delayed_10;
  b31_data_delayed_12 <= b31_data_delayed_11;
  b31_data_delayed_13 <= b31_data_delayed_12;
  b31_data_delayed_14 <= b31_data_delayed_13;
  b31_data_delayed_15 <= b31_data_delayed_14;
  b31_data_delayed_16 <= b31_data_delayed_15;
  b31_data_delayed_17 <= b31_data_delayed_16;
  b31_data_delayed_18 <= b31_data_delayed_17;
  b31_data_delayed_19 <= b31_data_delayed_18;
  b31_data_delayed_20 <= b31_data_delayed_19;
  b31_data_delayed_21 <= b31_data_delayed_20;
  b31_data_delayed_22 <= b31_data_delayed_21;
  b31_data_delayed_23 <= b31_data_delayed_22;
  b31_data_delayed_24 <= b31_data_delayed_23;
  b31_data_delayed_25 <= b31_data_delayed_24;
  b31_data_delayed_26 <= b31_data_delayed_25;
  b31_data_delayed_27 <= b31_data_delayed_26;
  b31_data_delayed_28 <= b31_data_delayed_27;
  b31_data_delayed_29 <= b31_data_delayed_28;
  b31_data_delayed_30 <= b31_data_delayed_29;
  b31_data_delayed_31 <= b31_data_delayed_30;
 
  end
end
endmodule


//////////////////////////////////////////////////////////////////////////
// Systolically connected PEs
//////////////////////////////////////////////////////////////////////////
module systolic_pe_matrix(
clk,
reset,
pe_reset,
start_mat_mul,
a0,
a1,
a2,
a3,
a4,
a5,
a6,
a7,
a8,
a9,
a10,
a11,
a12,
a13,
a14,
a15,
a16,
a17,
a18,
a19,
a20,
a21,
a22,
a23,
a24,
a25,
a26,
a27,
a28,
a29,
a30,
a31,
b0,
b1,
b2,
b3,
b4,
b5,
b6,
b7,
b8,
b9,
b10,
b11,
b12,
b13,
b14,
b15,
b16,
b17,
b18,
b19,
b20,
b21,
b22,
b23,
b24,
b25,
b26,
b27,
b28,
b29,
b30,
b31,
matrixC0_0,
matrixC0_1,
matrixC0_2,
matrixC0_3,
matrixC0_4,
matrixC0_5,
matrixC0_6,
matrixC0_7,
matrixC0_8,
matrixC0_9,
matrixC0_10,
matrixC0_11,
matrixC0_12,
matrixC0_13,
matrixC0_14,
matrixC0_15,
matrixC0_16,
matrixC0_17,
matrixC0_18,
matrixC0_19,
matrixC0_20,
matrixC0_21,
matrixC0_22,
matrixC0_23,
matrixC0_24,
matrixC0_25,
matrixC0_26,
matrixC0_27,
matrixC0_28,
matrixC0_29,
matrixC0_30,
matrixC0_31,
matrixC1_0,
matrixC1_1,
matrixC1_2,
matrixC1_3,
matrixC1_4,
matrixC1_5,
matrixC1_6,
matrixC1_7,
matrixC1_8,
matrixC1_9,
matrixC1_10,
matrixC1_11,
matrixC1_12,
matrixC1_13,
matrixC1_14,
matrixC1_15,
matrixC1_16,
matrixC1_17,
matrixC1_18,
matrixC1_19,
matrixC1_20,
matrixC1_21,
matrixC1_22,
matrixC1_23,
matrixC1_24,
matrixC1_25,
matrixC1_26,
matrixC1_27,
matrixC1_28,
matrixC1_29,
matrixC1_30,
matrixC1_31,
matrixC2_0,
matrixC2_1,
matrixC2_2,
matrixC2_3,
matrixC2_4,
matrixC2_5,
matrixC2_6,
matrixC2_7,
matrixC2_8,
matrixC2_9,
matrixC2_10,
matrixC2_11,
matrixC2_12,
matrixC2_13,
matrixC2_14,
matrixC2_15,
matrixC2_16,
matrixC2_17,
matrixC2_18,
matrixC2_19,
matrixC2_20,
matrixC2_21,
matrixC2_22,
matrixC2_23,
matrixC2_24,
matrixC2_25,
matrixC2_26,
matrixC2_27,
matrixC2_28,
matrixC2_29,
matrixC2_30,
matrixC2_31,
matrixC3_0,
matrixC3_1,
matrixC3_2,
matrixC3_3,
matrixC3_4,
matrixC3_5,
matrixC3_6,
matrixC3_7,
matrixC3_8,
matrixC3_9,
matrixC3_10,
matrixC3_11,
matrixC3_12,
matrixC3_13,
matrixC3_14,
matrixC3_15,
matrixC3_16,
matrixC3_17,
matrixC3_18,
matrixC3_19,
matrixC3_20,
matrixC3_21,
matrixC3_22,
matrixC3_23,
matrixC3_24,
matrixC3_25,
matrixC3_26,
matrixC3_27,
matrixC3_28,
matrixC3_29,
matrixC3_30,
matrixC3_31,
matrixC4_0,
matrixC4_1,
matrixC4_2,
matrixC4_3,
matrixC4_4,
matrixC4_5,
matrixC4_6,
matrixC4_7,
matrixC4_8,
matrixC4_9,
matrixC4_10,
matrixC4_11,
matrixC4_12,
matrixC4_13,
matrixC4_14,
matrixC4_15,
matrixC4_16,
matrixC4_17,
matrixC4_18,
matrixC4_19,
matrixC4_20,
matrixC4_21,
matrixC4_22,
matrixC4_23,
matrixC4_24,
matrixC4_25,
matrixC4_26,
matrixC4_27,
matrixC4_28,
matrixC4_29,
matrixC4_30,
matrixC4_31,
matrixC5_0,
matrixC5_1,
matrixC5_2,
matrixC5_3,
matrixC5_4,
matrixC5_5,
matrixC5_6,
matrixC5_7,
matrixC5_8,
matrixC5_9,
matrixC5_10,
matrixC5_11,
matrixC5_12,
matrixC5_13,
matrixC5_14,
matrixC5_15,
matrixC5_16,
matrixC5_17,
matrixC5_18,
matrixC5_19,
matrixC5_20,
matrixC5_21,
matrixC5_22,
matrixC5_23,
matrixC5_24,
matrixC5_25,
matrixC5_26,
matrixC5_27,
matrixC5_28,
matrixC5_29,
matrixC5_30,
matrixC5_31,
matrixC6_0,
matrixC6_1,
matrixC6_2,
matrixC6_3,
matrixC6_4,
matrixC6_5,
matrixC6_6,
matrixC6_7,
matrixC6_8,
matrixC6_9,
matrixC6_10,
matrixC6_11,
matrixC6_12,
matrixC6_13,
matrixC6_14,
matrixC6_15,
matrixC6_16,
matrixC6_17,
matrixC6_18,
matrixC6_19,
matrixC6_20,
matrixC6_21,
matrixC6_22,
matrixC6_23,
matrixC6_24,
matrixC6_25,
matrixC6_26,
matrixC6_27,
matrixC6_28,
matrixC6_29,
matrixC6_30,
matrixC6_31,
matrixC7_0,
matrixC7_1,
matrixC7_2,
matrixC7_3,
matrixC7_4,
matrixC7_5,
matrixC7_6,
matrixC7_7,
matrixC7_8,
matrixC7_9,
matrixC7_10,
matrixC7_11,
matrixC7_12,
matrixC7_13,
matrixC7_14,
matrixC7_15,
matrixC7_16,
matrixC7_17,
matrixC7_18,
matrixC7_19,
matrixC7_20,
matrixC7_21,
matrixC7_22,
matrixC7_23,
matrixC7_24,
matrixC7_25,
matrixC7_26,
matrixC7_27,
matrixC7_28,
matrixC7_29,
matrixC7_30,
matrixC7_31,
matrixC8_0,
matrixC8_1,
matrixC8_2,
matrixC8_3,
matrixC8_4,
matrixC8_5,
matrixC8_6,
matrixC8_7,
matrixC8_8,
matrixC8_9,
matrixC8_10,
matrixC8_11,
matrixC8_12,
matrixC8_13,
matrixC8_14,
matrixC8_15,
matrixC8_16,
matrixC8_17,
matrixC8_18,
matrixC8_19,
matrixC8_20,
matrixC8_21,
matrixC8_22,
matrixC8_23,
matrixC8_24,
matrixC8_25,
matrixC8_26,
matrixC8_27,
matrixC8_28,
matrixC8_29,
matrixC8_30,
matrixC8_31,
matrixC9_0,
matrixC9_1,
matrixC9_2,
matrixC9_3,
matrixC9_4,
matrixC9_5,
matrixC9_6,
matrixC9_7,
matrixC9_8,
matrixC9_9,
matrixC9_10,
matrixC9_11,
matrixC9_12,
matrixC9_13,
matrixC9_14,
matrixC9_15,
matrixC9_16,
matrixC9_17,
matrixC9_18,
matrixC9_19,
matrixC9_20,
matrixC9_21,
matrixC9_22,
matrixC9_23,
matrixC9_24,
matrixC9_25,
matrixC9_26,
matrixC9_27,
matrixC9_28,
matrixC9_29,
matrixC9_30,
matrixC9_31,
matrixC10_0,
matrixC10_1,
matrixC10_2,
matrixC10_3,
matrixC10_4,
matrixC10_5,
matrixC10_6,
matrixC10_7,
matrixC10_8,
matrixC10_9,
matrixC10_10,
matrixC10_11,
matrixC10_12,
matrixC10_13,
matrixC10_14,
matrixC10_15,
matrixC10_16,
matrixC10_17,
matrixC10_18,
matrixC10_19,
matrixC10_20,
matrixC10_21,
matrixC10_22,
matrixC10_23,
matrixC10_24,
matrixC10_25,
matrixC10_26,
matrixC10_27,
matrixC10_28,
matrixC10_29,
matrixC10_30,
matrixC10_31,
matrixC11_0,
matrixC11_1,
matrixC11_2,
matrixC11_3,
matrixC11_4,
matrixC11_5,
matrixC11_6,
matrixC11_7,
matrixC11_8,
matrixC11_9,
matrixC11_10,
matrixC11_11,
matrixC11_12,
matrixC11_13,
matrixC11_14,
matrixC11_15,
matrixC11_16,
matrixC11_17,
matrixC11_18,
matrixC11_19,
matrixC11_20,
matrixC11_21,
matrixC11_22,
matrixC11_23,
matrixC11_24,
matrixC11_25,
matrixC11_26,
matrixC11_27,
matrixC11_28,
matrixC11_29,
matrixC11_30,
matrixC11_31,
matrixC12_0,
matrixC12_1,
matrixC12_2,
matrixC12_3,
matrixC12_4,
matrixC12_5,
matrixC12_6,
matrixC12_7,
matrixC12_8,
matrixC12_9,
matrixC12_10,
matrixC12_11,
matrixC12_12,
matrixC12_13,
matrixC12_14,
matrixC12_15,
matrixC12_16,
matrixC12_17,
matrixC12_18,
matrixC12_19,
matrixC12_20,
matrixC12_21,
matrixC12_22,
matrixC12_23,
matrixC12_24,
matrixC12_25,
matrixC12_26,
matrixC12_27,
matrixC12_28,
matrixC12_29,
matrixC12_30,
matrixC12_31,
matrixC13_0,
matrixC13_1,
matrixC13_2,
matrixC13_3,
matrixC13_4,
matrixC13_5,
matrixC13_6,
matrixC13_7,
matrixC13_8,
matrixC13_9,
matrixC13_10,
matrixC13_11,
matrixC13_12,
matrixC13_13,
matrixC13_14,
matrixC13_15,
matrixC13_16,
matrixC13_17,
matrixC13_18,
matrixC13_19,
matrixC13_20,
matrixC13_21,
matrixC13_22,
matrixC13_23,
matrixC13_24,
matrixC13_25,
matrixC13_26,
matrixC13_27,
matrixC13_28,
matrixC13_29,
matrixC13_30,
matrixC13_31,
matrixC14_0,
matrixC14_1,
matrixC14_2,
matrixC14_3,
matrixC14_4,
matrixC14_5,
matrixC14_6,
matrixC14_7,
matrixC14_8,
matrixC14_9,
matrixC14_10,
matrixC14_11,
matrixC14_12,
matrixC14_13,
matrixC14_14,
matrixC14_15,
matrixC14_16,
matrixC14_17,
matrixC14_18,
matrixC14_19,
matrixC14_20,
matrixC14_21,
matrixC14_22,
matrixC14_23,
matrixC14_24,
matrixC14_25,
matrixC14_26,
matrixC14_27,
matrixC14_28,
matrixC14_29,
matrixC14_30,
matrixC14_31,
matrixC15_0,
matrixC15_1,
matrixC15_2,
matrixC15_3,
matrixC15_4,
matrixC15_5,
matrixC15_6,
matrixC15_7,
matrixC15_8,
matrixC15_9,
matrixC15_10,
matrixC15_11,
matrixC15_12,
matrixC15_13,
matrixC15_14,
matrixC15_15,
matrixC15_16,
matrixC15_17,
matrixC15_18,
matrixC15_19,
matrixC15_20,
matrixC15_21,
matrixC15_22,
matrixC15_23,
matrixC15_24,
matrixC15_25,
matrixC15_26,
matrixC15_27,
matrixC15_28,
matrixC15_29,
matrixC15_30,
matrixC15_31,
matrixC16_0,
matrixC16_1,
matrixC16_2,
matrixC16_3,
matrixC16_4,
matrixC16_5,
matrixC16_6,
matrixC16_7,
matrixC16_8,
matrixC16_9,
matrixC16_10,
matrixC16_11,
matrixC16_12,
matrixC16_13,
matrixC16_14,
matrixC16_15,
matrixC16_16,
matrixC16_17,
matrixC16_18,
matrixC16_19,
matrixC16_20,
matrixC16_21,
matrixC16_22,
matrixC16_23,
matrixC16_24,
matrixC16_25,
matrixC16_26,
matrixC16_27,
matrixC16_28,
matrixC16_29,
matrixC16_30,
matrixC16_31,
matrixC17_0,
matrixC17_1,
matrixC17_2,
matrixC17_3,
matrixC17_4,
matrixC17_5,
matrixC17_6,
matrixC17_7,
matrixC17_8,
matrixC17_9,
matrixC17_10,
matrixC17_11,
matrixC17_12,
matrixC17_13,
matrixC17_14,
matrixC17_15,
matrixC17_16,
matrixC17_17,
matrixC17_18,
matrixC17_19,
matrixC17_20,
matrixC17_21,
matrixC17_22,
matrixC17_23,
matrixC17_24,
matrixC17_25,
matrixC17_26,
matrixC17_27,
matrixC17_28,
matrixC17_29,
matrixC17_30,
matrixC17_31,
matrixC18_0,
matrixC18_1,
matrixC18_2,
matrixC18_3,
matrixC18_4,
matrixC18_5,
matrixC18_6,
matrixC18_7,
matrixC18_8,
matrixC18_9,
matrixC18_10,
matrixC18_11,
matrixC18_12,
matrixC18_13,
matrixC18_14,
matrixC18_15,
matrixC18_16,
matrixC18_17,
matrixC18_18,
matrixC18_19,
matrixC18_20,
matrixC18_21,
matrixC18_22,
matrixC18_23,
matrixC18_24,
matrixC18_25,
matrixC18_26,
matrixC18_27,
matrixC18_28,
matrixC18_29,
matrixC18_30,
matrixC18_31,
matrixC19_0,
matrixC19_1,
matrixC19_2,
matrixC19_3,
matrixC19_4,
matrixC19_5,
matrixC19_6,
matrixC19_7,
matrixC19_8,
matrixC19_9,
matrixC19_10,
matrixC19_11,
matrixC19_12,
matrixC19_13,
matrixC19_14,
matrixC19_15,
matrixC19_16,
matrixC19_17,
matrixC19_18,
matrixC19_19,
matrixC19_20,
matrixC19_21,
matrixC19_22,
matrixC19_23,
matrixC19_24,
matrixC19_25,
matrixC19_26,
matrixC19_27,
matrixC19_28,
matrixC19_29,
matrixC19_30,
matrixC19_31,
matrixC20_0,
matrixC20_1,
matrixC20_2,
matrixC20_3,
matrixC20_4,
matrixC20_5,
matrixC20_6,
matrixC20_7,
matrixC20_8,
matrixC20_9,
matrixC20_10,
matrixC20_11,
matrixC20_12,
matrixC20_13,
matrixC20_14,
matrixC20_15,
matrixC20_16,
matrixC20_17,
matrixC20_18,
matrixC20_19,
matrixC20_20,
matrixC20_21,
matrixC20_22,
matrixC20_23,
matrixC20_24,
matrixC20_25,
matrixC20_26,
matrixC20_27,
matrixC20_28,
matrixC20_29,
matrixC20_30,
matrixC20_31,
matrixC21_0,
matrixC21_1,
matrixC21_2,
matrixC21_3,
matrixC21_4,
matrixC21_5,
matrixC21_6,
matrixC21_7,
matrixC21_8,
matrixC21_9,
matrixC21_10,
matrixC21_11,
matrixC21_12,
matrixC21_13,
matrixC21_14,
matrixC21_15,
matrixC21_16,
matrixC21_17,
matrixC21_18,
matrixC21_19,
matrixC21_20,
matrixC21_21,
matrixC21_22,
matrixC21_23,
matrixC21_24,
matrixC21_25,
matrixC21_26,
matrixC21_27,
matrixC21_28,
matrixC21_29,
matrixC21_30,
matrixC21_31,
matrixC22_0,
matrixC22_1,
matrixC22_2,
matrixC22_3,
matrixC22_4,
matrixC22_5,
matrixC22_6,
matrixC22_7,
matrixC22_8,
matrixC22_9,
matrixC22_10,
matrixC22_11,
matrixC22_12,
matrixC22_13,
matrixC22_14,
matrixC22_15,
matrixC22_16,
matrixC22_17,
matrixC22_18,
matrixC22_19,
matrixC22_20,
matrixC22_21,
matrixC22_22,
matrixC22_23,
matrixC22_24,
matrixC22_25,
matrixC22_26,
matrixC22_27,
matrixC22_28,
matrixC22_29,
matrixC22_30,
matrixC22_31,
matrixC23_0,
matrixC23_1,
matrixC23_2,
matrixC23_3,
matrixC23_4,
matrixC23_5,
matrixC23_6,
matrixC23_7,
matrixC23_8,
matrixC23_9,
matrixC23_10,
matrixC23_11,
matrixC23_12,
matrixC23_13,
matrixC23_14,
matrixC23_15,
matrixC23_16,
matrixC23_17,
matrixC23_18,
matrixC23_19,
matrixC23_20,
matrixC23_21,
matrixC23_22,
matrixC23_23,
matrixC23_24,
matrixC23_25,
matrixC23_26,
matrixC23_27,
matrixC23_28,
matrixC23_29,
matrixC23_30,
matrixC23_31,
matrixC24_0,
matrixC24_1,
matrixC24_2,
matrixC24_3,
matrixC24_4,
matrixC24_5,
matrixC24_6,
matrixC24_7,
matrixC24_8,
matrixC24_9,
matrixC24_10,
matrixC24_11,
matrixC24_12,
matrixC24_13,
matrixC24_14,
matrixC24_15,
matrixC24_16,
matrixC24_17,
matrixC24_18,
matrixC24_19,
matrixC24_20,
matrixC24_21,
matrixC24_22,
matrixC24_23,
matrixC24_24,
matrixC24_25,
matrixC24_26,
matrixC24_27,
matrixC24_28,
matrixC24_29,
matrixC24_30,
matrixC24_31,
matrixC25_0,
matrixC25_1,
matrixC25_2,
matrixC25_3,
matrixC25_4,
matrixC25_5,
matrixC25_6,
matrixC25_7,
matrixC25_8,
matrixC25_9,
matrixC25_10,
matrixC25_11,
matrixC25_12,
matrixC25_13,
matrixC25_14,
matrixC25_15,
matrixC25_16,
matrixC25_17,
matrixC25_18,
matrixC25_19,
matrixC25_20,
matrixC25_21,
matrixC25_22,
matrixC25_23,
matrixC25_24,
matrixC25_25,
matrixC25_26,
matrixC25_27,
matrixC25_28,
matrixC25_29,
matrixC25_30,
matrixC25_31,
matrixC26_0,
matrixC26_1,
matrixC26_2,
matrixC26_3,
matrixC26_4,
matrixC26_5,
matrixC26_6,
matrixC26_7,
matrixC26_8,
matrixC26_9,
matrixC26_10,
matrixC26_11,
matrixC26_12,
matrixC26_13,
matrixC26_14,
matrixC26_15,
matrixC26_16,
matrixC26_17,
matrixC26_18,
matrixC26_19,
matrixC26_20,
matrixC26_21,
matrixC26_22,
matrixC26_23,
matrixC26_24,
matrixC26_25,
matrixC26_26,
matrixC26_27,
matrixC26_28,
matrixC26_29,
matrixC26_30,
matrixC26_31,
matrixC27_0,
matrixC27_1,
matrixC27_2,
matrixC27_3,
matrixC27_4,
matrixC27_5,
matrixC27_6,
matrixC27_7,
matrixC27_8,
matrixC27_9,
matrixC27_10,
matrixC27_11,
matrixC27_12,
matrixC27_13,
matrixC27_14,
matrixC27_15,
matrixC27_16,
matrixC27_17,
matrixC27_18,
matrixC27_19,
matrixC27_20,
matrixC27_21,
matrixC27_22,
matrixC27_23,
matrixC27_24,
matrixC27_25,
matrixC27_26,
matrixC27_27,
matrixC27_28,
matrixC27_29,
matrixC27_30,
matrixC27_31,
matrixC28_0,
matrixC28_1,
matrixC28_2,
matrixC28_3,
matrixC28_4,
matrixC28_5,
matrixC28_6,
matrixC28_7,
matrixC28_8,
matrixC28_9,
matrixC28_10,
matrixC28_11,
matrixC28_12,
matrixC28_13,
matrixC28_14,
matrixC28_15,
matrixC28_16,
matrixC28_17,
matrixC28_18,
matrixC28_19,
matrixC28_20,
matrixC28_21,
matrixC28_22,
matrixC28_23,
matrixC28_24,
matrixC28_25,
matrixC28_26,
matrixC28_27,
matrixC28_28,
matrixC28_29,
matrixC28_30,
matrixC28_31,
matrixC29_0,
matrixC29_1,
matrixC29_2,
matrixC29_3,
matrixC29_4,
matrixC29_5,
matrixC29_6,
matrixC29_7,
matrixC29_8,
matrixC29_9,
matrixC29_10,
matrixC29_11,
matrixC29_12,
matrixC29_13,
matrixC29_14,
matrixC29_15,
matrixC29_16,
matrixC29_17,
matrixC29_18,
matrixC29_19,
matrixC29_20,
matrixC29_21,
matrixC29_22,
matrixC29_23,
matrixC29_24,
matrixC29_25,
matrixC29_26,
matrixC29_27,
matrixC29_28,
matrixC29_29,
matrixC29_30,
matrixC29_31,
matrixC30_0,
matrixC30_1,
matrixC30_2,
matrixC30_3,
matrixC30_4,
matrixC30_5,
matrixC30_6,
matrixC30_7,
matrixC30_8,
matrixC30_9,
matrixC30_10,
matrixC30_11,
matrixC30_12,
matrixC30_13,
matrixC30_14,
matrixC30_15,
matrixC30_16,
matrixC30_17,
matrixC30_18,
matrixC30_19,
matrixC30_20,
matrixC30_21,
matrixC30_22,
matrixC30_23,
matrixC30_24,
matrixC30_25,
matrixC30_26,
matrixC30_27,
matrixC30_28,
matrixC30_29,
matrixC30_30,
matrixC30_31,
matrixC31_0,
matrixC31_1,
matrixC31_2,
matrixC31_3,
matrixC31_4,
matrixC31_5,
matrixC31_6,
matrixC31_7,
matrixC31_8,
matrixC31_9,
matrixC31_10,
matrixC31_11,
matrixC31_12,
matrixC31_13,
matrixC31_14,
matrixC31_15,
matrixC31_16,
matrixC31_17,
matrixC31_18,
matrixC31_19,
matrixC31_20,
matrixC31_21,
matrixC31_22,
matrixC31_23,
matrixC31_24,
matrixC31_25,
matrixC31_26,
matrixC31_27,
matrixC31_28,
matrixC31_29,
matrixC31_30,
matrixC31_31,

a_data_out,
b_data_out
);

input clk;
input reset;
input pe_reset;
input start_mat_mul;
input [`DWIDTH-1:0] a0;
input [`DWIDTH-1:0] a1;
input [`DWIDTH-1:0] a2;
input [`DWIDTH-1:0] a3;
input [`DWIDTH-1:0] a4;
input [`DWIDTH-1:0] a5;
input [`DWIDTH-1:0] a6;
input [`DWIDTH-1:0] a7;
input [`DWIDTH-1:0] a8;
input [`DWIDTH-1:0] a9;
input [`DWIDTH-1:0] a10;
input [`DWIDTH-1:0] a11;
input [`DWIDTH-1:0] a12;
input [`DWIDTH-1:0] a13;
input [`DWIDTH-1:0] a14;
input [`DWIDTH-1:0] a15;
input [`DWIDTH-1:0] a16;
input [`DWIDTH-1:0] a17;
input [`DWIDTH-1:0] a18;
input [`DWIDTH-1:0] a19;
input [`DWIDTH-1:0] a20;
input [`DWIDTH-1:0] a21;
input [`DWIDTH-1:0] a22;
input [`DWIDTH-1:0] a23;
input [`DWIDTH-1:0] a24;
input [`DWIDTH-1:0] a25;
input [`DWIDTH-1:0] a26;
input [`DWIDTH-1:0] a27;
input [`DWIDTH-1:0] a28;
input [`DWIDTH-1:0] a29;
input [`DWIDTH-1:0] a30;
input [`DWIDTH-1:0] a31;
input [`DWIDTH-1:0] b0;
input [`DWIDTH-1:0] b1;
input [`DWIDTH-1:0] b2;
input [`DWIDTH-1:0] b3;
input [`DWIDTH-1:0] b4;
input [`DWIDTH-1:0] b5;
input [`DWIDTH-1:0] b6;
input [`DWIDTH-1:0] b7;
input [`DWIDTH-1:0] b8;
input [`DWIDTH-1:0] b9;
input [`DWIDTH-1:0] b10;
input [`DWIDTH-1:0] b11;
input [`DWIDTH-1:0] b12;
input [`DWIDTH-1:0] b13;
input [`DWIDTH-1:0] b14;
input [`DWIDTH-1:0] b15;
input [`DWIDTH-1:0] b16;
input [`DWIDTH-1:0] b17;
input [`DWIDTH-1:0] b18;
input [`DWIDTH-1:0] b19;
input [`DWIDTH-1:0] b20;
input [`DWIDTH-1:0] b21;
input [`DWIDTH-1:0] b22;
input [`DWIDTH-1:0] b23;
input [`DWIDTH-1:0] b24;
input [`DWIDTH-1:0] b25;
input [`DWIDTH-1:0] b26;
input [`DWIDTH-1:0] b27;
input [`DWIDTH-1:0] b28;
input [`DWIDTH-1:0] b29;
input [`DWIDTH-1:0] b30;
input [`DWIDTH-1:0] b31;
output [`DWIDTH-1:0] matrixC0_0;
output [`DWIDTH-1:0] matrixC0_1;
output [`DWIDTH-1:0] matrixC0_2;
output [`DWIDTH-1:0] matrixC0_3;
output [`DWIDTH-1:0] matrixC0_4;
output [`DWIDTH-1:0] matrixC0_5;
output [`DWIDTH-1:0] matrixC0_6;
output [`DWIDTH-1:0] matrixC0_7;
output [`DWIDTH-1:0] matrixC0_8;
output [`DWIDTH-1:0] matrixC0_9;
output [`DWIDTH-1:0] matrixC0_10;
output [`DWIDTH-1:0] matrixC0_11;
output [`DWIDTH-1:0] matrixC0_12;
output [`DWIDTH-1:0] matrixC0_13;
output [`DWIDTH-1:0] matrixC0_14;
output [`DWIDTH-1:0] matrixC0_15;
output [`DWIDTH-1:0] matrixC0_16;
output [`DWIDTH-1:0] matrixC0_17;
output [`DWIDTH-1:0] matrixC0_18;
output [`DWIDTH-1:0] matrixC0_19;
output [`DWIDTH-1:0] matrixC0_20;
output [`DWIDTH-1:0] matrixC0_21;
output [`DWIDTH-1:0] matrixC0_22;
output [`DWIDTH-1:0] matrixC0_23;
output [`DWIDTH-1:0] matrixC0_24;
output [`DWIDTH-1:0] matrixC0_25;
output [`DWIDTH-1:0] matrixC0_26;
output [`DWIDTH-1:0] matrixC0_27;
output [`DWIDTH-1:0] matrixC0_28;
output [`DWIDTH-1:0] matrixC0_29;
output [`DWIDTH-1:0] matrixC0_30;
output [`DWIDTH-1:0] matrixC0_31;
output [`DWIDTH-1:0] matrixC1_0;
output [`DWIDTH-1:0] matrixC1_1;
output [`DWIDTH-1:0] matrixC1_2;
output [`DWIDTH-1:0] matrixC1_3;
output [`DWIDTH-1:0] matrixC1_4;
output [`DWIDTH-1:0] matrixC1_5;
output [`DWIDTH-1:0] matrixC1_6;
output [`DWIDTH-1:0] matrixC1_7;
output [`DWIDTH-1:0] matrixC1_8;
output [`DWIDTH-1:0] matrixC1_9;
output [`DWIDTH-1:0] matrixC1_10;
output [`DWIDTH-1:0] matrixC1_11;
output [`DWIDTH-1:0] matrixC1_12;
output [`DWIDTH-1:0] matrixC1_13;
output [`DWIDTH-1:0] matrixC1_14;
output [`DWIDTH-1:0] matrixC1_15;
output [`DWIDTH-1:0] matrixC1_16;
output [`DWIDTH-1:0] matrixC1_17;
output [`DWIDTH-1:0] matrixC1_18;
output [`DWIDTH-1:0] matrixC1_19;
output [`DWIDTH-1:0] matrixC1_20;
output [`DWIDTH-1:0] matrixC1_21;
output [`DWIDTH-1:0] matrixC1_22;
output [`DWIDTH-1:0] matrixC1_23;
output [`DWIDTH-1:0] matrixC1_24;
output [`DWIDTH-1:0] matrixC1_25;
output [`DWIDTH-1:0] matrixC1_26;
output [`DWIDTH-1:0] matrixC1_27;
output [`DWIDTH-1:0] matrixC1_28;
output [`DWIDTH-1:0] matrixC1_29;
output [`DWIDTH-1:0] matrixC1_30;
output [`DWIDTH-1:0] matrixC1_31;
output [`DWIDTH-1:0] matrixC2_0;
output [`DWIDTH-1:0] matrixC2_1;
output [`DWIDTH-1:0] matrixC2_2;
output [`DWIDTH-1:0] matrixC2_3;
output [`DWIDTH-1:0] matrixC2_4;
output [`DWIDTH-1:0] matrixC2_5;
output [`DWIDTH-1:0] matrixC2_6;
output [`DWIDTH-1:0] matrixC2_7;
output [`DWIDTH-1:0] matrixC2_8;
output [`DWIDTH-1:0] matrixC2_9;
output [`DWIDTH-1:0] matrixC2_10;
output [`DWIDTH-1:0] matrixC2_11;
output [`DWIDTH-1:0] matrixC2_12;
output [`DWIDTH-1:0] matrixC2_13;
output [`DWIDTH-1:0] matrixC2_14;
output [`DWIDTH-1:0] matrixC2_15;
output [`DWIDTH-1:0] matrixC2_16;
output [`DWIDTH-1:0] matrixC2_17;
output [`DWIDTH-1:0] matrixC2_18;
output [`DWIDTH-1:0] matrixC2_19;
output [`DWIDTH-1:0] matrixC2_20;
output [`DWIDTH-1:0] matrixC2_21;
output [`DWIDTH-1:0] matrixC2_22;
output [`DWIDTH-1:0] matrixC2_23;
output [`DWIDTH-1:0] matrixC2_24;
output [`DWIDTH-1:0] matrixC2_25;
output [`DWIDTH-1:0] matrixC2_26;
output [`DWIDTH-1:0] matrixC2_27;
output [`DWIDTH-1:0] matrixC2_28;
output [`DWIDTH-1:0] matrixC2_29;
output [`DWIDTH-1:0] matrixC2_30;
output [`DWIDTH-1:0] matrixC2_31;
output [`DWIDTH-1:0] matrixC3_0;
output [`DWIDTH-1:0] matrixC3_1;
output [`DWIDTH-1:0] matrixC3_2;
output [`DWIDTH-1:0] matrixC3_3;
output [`DWIDTH-1:0] matrixC3_4;
output [`DWIDTH-1:0] matrixC3_5;
output [`DWIDTH-1:0] matrixC3_6;
output [`DWIDTH-1:0] matrixC3_7;
output [`DWIDTH-1:0] matrixC3_8;
output [`DWIDTH-1:0] matrixC3_9;
output [`DWIDTH-1:0] matrixC3_10;
output [`DWIDTH-1:0] matrixC3_11;
output [`DWIDTH-1:0] matrixC3_12;
output [`DWIDTH-1:0] matrixC3_13;
output [`DWIDTH-1:0] matrixC3_14;
output [`DWIDTH-1:0] matrixC3_15;
output [`DWIDTH-1:0] matrixC3_16;
output [`DWIDTH-1:0] matrixC3_17;
output [`DWIDTH-1:0] matrixC3_18;
output [`DWIDTH-1:0] matrixC3_19;
output [`DWIDTH-1:0] matrixC3_20;
output [`DWIDTH-1:0] matrixC3_21;
output [`DWIDTH-1:0] matrixC3_22;
output [`DWIDTH-1:0] matrixC3_23;
output [`DWIDTH-1:0] matrixC3_24;
output [`DWIDTH-1:0] matrixC3_25;
output [`DWIDTH-1:0] matrixC3_26;
output [`DWIDTH-1:0] matrixC3_27;
output [`DWIDTH-1:0] matrixC3_28;
output [`DWIDTH-1:0] matrixC3_29;
output [`DWIDTH-1:0] matrixC3_30;
output [`DWIDTH-1:0] matrixC3_31;
output [`DWIDTH-1:0] matrixC4_0;
output [`DWIDTH-1:0] matrixC4_1;
output [`DWIDTH-1:0] matrixC4_2;
output [`DWIDTH-1:0] matrixC4_3;
output [`DWIDTH-1:0] matrixC4_4;
output [`DWIDTH-1:0] matrixC4_5;
output [`DWIDTH-1:0] matrixC4_6;
output [`DWIDTH-1:0] matrixC4_7;
output [`DWIDTH-1:0] matrixC4_8;
output [`DWIDTH-1:0] matrixC4_9;
output [`DWIDTH-1:0] matrixC4_10;
output [`DWIDTH-1:0] matrixC4_11;
output [`DWIDTH-1:0] matrixC4_12;
output [`DWIDTH-1:0] matrixC4_13;
output [`DWIDTH-1:0] matrixC4_14;
output [`DWIDTH-1:0] matrixC4_15;
output [`DWIDTH-1:0] matrixC4_16;
output [`DWIDTH-1:0] matrixC4_17;
output [`DWIDTH-1:0] matrixC4_18;
output [`DWIDTH-1:0] matrixC4_19;
output [`DWIDTH-1:0] matrixC4_20;
output [`DWIDTH-1:0] matrixC4_21;
output [`DWIDTH-1:0] matrixC4_22;
output [`DWIDTH-1:0] matrixC4_23;
output [`DWIDTH-1:0] matrixC4_24;
output [`DWIDTH-1:0] matrixC4_25;
output [`DWIDTH-1:0] matrixC4_26;
output [`DWIDTH-1:0] matrixC4_27;
output [`DWIDTH-1:0] matrixC4_28;
output [`DWIDTH-1:0] matrixC4_29;
output [`DWIDTH-1:0] matrixC4_30;
output [`DWIDTH-1:0] matrixC4_31;
output [`DWIDTH-1:0] matrixC5_0;
output [`DWIDTH-1:0] matrixC5_1;
output [`DWIDTH-1:0] matrixC5_2;
output [`DWIDTH-1:0] matrixC5_3;
output [`DWIDTH-1:0] matrixC5_4;
output [`DWIDTH-1:0] matrixC5_5;
output [`DWIDTH-1:0] matrixC5_6;
output [`DWIDTH-1:0] matrixC5_7;
output [`DWIDTH-1:0] matrixC5_8;
output [`DWIDTH-1:0] matrixC5_9;
output [`DWIDTH-1:0] matrixC5_10;
output [`DWIDTH-1:0] matrixC5_11;
output [`DWIDTH-1:0] matrixC5_12;
output [`DWIDTH-1:0] matrixC5_13;
output [`DWIDTH-1:0] matrixC5_14;
output [`DWIDTH-1:0] matrixC5_15;
output [`DWIDTH-1:0] matrixC5_16;
output [`DWIDTH-1:0] matrixC5_17;
output [`DWIDTH-1:0] matrixC5_18;
output [`DWIDTH-1:0] matrixC5_19;
output [`DWIDTH-1:0] matrixC5_20;
output [`DWIDTH-1:0] matrixC5_21;
output [`DWIDTH-1:0] matrixC5_22;
output [`DWIDTH-1:0] matrixC5_23;
output [`DWIDTH-1:0] matrixC5_24;
output [`DWIDTH-1:0] matrixC5_25;
output [`DWIDTH-1:0] matrixC5_26;
output [`DWIDTH-1:0] matrixC5_27;
output [`DWIDTH-1:0] matrixC5_28;
output [`DWIDTH-1:0] matrixC5_29;
output [`DWIDTH-1:0] matrixC5_30;
output [`DWIDTH-1:0] matrixC5_31;
output [`DWIDTH-1:0] matrixC6_0;
output [`DWIDTH-1:0] matrixC6_1;
output [`DWIDTH-1:0] matrixC6_2;
output [`DWIDTH-1:0] matrixC6_3;
output [`DWIDTH-1:0] matrixC6_4;
output [`DWIDTH-1:0] matrixC6_5;
output [`DWIDTH-1:0] matrixC6_6;
output [`DWIDTH-1:0] matrixC6_7;
output [`DWIDTH-1:0] matrixC6_8;
output [`DWIDTH-1:0] matrixC6_9;
output [`DWIDTH-1:0] matrixC6_10;
output [`DWIDTH-1:0] matrixC6_11;
output [`DWIDTH-1:0] matrixC6_12;
output [`DWIDTH-1:0] matrixC6_13;
output [`DWIDTH-1:0] matrixC6_14;
output [`DWIDTH-1:0] matrixC6_15;
output [`DWIDTH-1:0] matrixC6_16;
output [`DWIDTH-1:0] matrixC6_17;
output [`DWIDTH-1:0] matrixC6_18;
output [`DWIDTH-1:0] matrixC6_19;
output [`DWIDTH-1:0] matrixC6_20;
output [`DWIDTH-1:0] matrixC6_21;
output [`DWIDTH-1:0] matrixC6_22;
output [`DWIDTH-1:0] matrixC6_23;
output [`DWIDTH-1:0] matrixC6_24;
output [`DWIDTH-1:0] matrixC6_25;
output [`DWIDTH-1:0] matrixC6_26;
output [`DWIDTH-1:0] matrixC6_27;
output [`DWIDTH-1:0] matrixC6_28;
output [`DWIDTH-1:0] matrixC6_29;
output [`DWIDTH-1:0] matrixC6_30;
output [`DWIDTH-1:0] matrixC6_31;
output [`DWIDTH-1:0] matrixC7_0;
output [`DWIDTH-1:0] matrixC7_1;
output [`DWIDTH-1:0] matrixC7_2;
output [`DWIDTH-1:0] matrixC7_3;
output [`DWIDTH-1:0] matrixC7_4;
output [`DWIDTH-1:0] matrixC7_5;
output [`DWIDTH-1:0] matrixC7_6;
output [`DWIDTH-1:0] matrixC7_7;
output [`DWIDTH-1:0] matrixC7_8;
output [`DWIDTH-1:0] matrixC7_9;
output [`DWIDTH-1:0] matrixC7_10;
output [`DWIDTH-1:0] matrixC7_11;
output [`DWIDTH-1:0] matrixC7_12;
output [`DWIDTH-1:0] matrixC7_13;
output [`DWIDTH-1:0] matrixC7_14;
output [`DWIDTH-1:0] matrixC7_15;
output [`DWIDTH-1:0] matrixC7_16;
output [`DWIDTH-1:0] matrixC7_17;
output [`DWIDTH-1:0] matrixC7_18;
output [`DWIDTH-1:0] matrixC7_19;
output [`DWIDTH-1:0] matrixC7_20;
output [`DWIDTH-1:0] matrixC7_21;
output [`DWIDTH-1:0] matrixC7_22;
output [`DWIDTH-1:0] matrixC7_23;
output [`DWIDTH-1:0] matrixC7_24;
output [`DWIDTH-1:0] matrixC7_25;
output [`DWIDTH-1:0] matrixC7_26;
output [`DWIDTH-1:0] matrixC7_27;
output [`DWIDTH-1:0] matrixC7_28;
output [`DWIDTH-1:0] matrixC7_29;
output [`DWIDTH-1:0] matrixC7_30;
output [`DWIDTH-1:0] matrixC7_31;
output [`DWIDTH-1:0] matrixC8_0;
output [`DWIDTH-1:0] matrixC8_1;
output [`DWIDTH-1:0] matrixC8_2;
output [`DWIDTH-1:0] matrixC8_3;
output [`DWIDTH-1:0] matrixC8_4;
output [`DWIDTH-1:0] matrixC8_5;
output [`DWIDTH-1:0] matrixC8_6;
output [`DWIDTH-1:0] matrixC8_7;
output [`DWIDTH-1:0] matrixC8_8;
output [`DWIDTH-1:0] matrixC8_9;
output [`DWIDTH-1:0] matrixC8_10;
output [`DWIDTH-1:0] matrixC8_11;
output [`DWIDTH-1:0] matrixC8_12;
output [`DWIDTH-1:0] matrixC8_13;
output [`DWIDTH-1:0] matrixC8_14;
output [`DWIDTH-1:0] matrixC8_15;
output [`DWIDTH-1:0] matrixC8_16;
output [`DWIDTH-1:0] matrixC8_17;
output [`DWIDTH-1:0] matrixC8_18;
output [`DWIDTH-1:0] matrixC8_19;
output [`DWIDTH-1:0] matrixC8_20;
output [`DWIDTH-1:0] matrixC8_21;
output [`DWIDTH-1:0] matrixC8_22;
output [`DWIDTH-1:0] matrixC8_23;
output [`DWIDTH-1:0] matrixC8_24;
output [`DWIDTH-1:0] matrixC8_25;
output [`DWIDTH-1:0] matrixC8_26;
output [`DWIDTH-1:0] matrixC8_27;
output [`DWIDTH-1:0] matrixC8_28;
output [`DWIDTH-1:0] matrixC8_29;
output [`DWIDTH-1:0] matrixC8_30;
output [`DWIDTH-1:0] matrixC8_31;
output [`DWIDTH-1:0] matrixC9_0;
output [`DWIDTH-1:0] matrixC9_1;
output [`DWIDTH-1:0] matrixC9_2;
output [`DWIDTH-1:0] matrixC9_3;
output [`DWIDTH-1:0] matrixC9_4;
output [`DWIDTH-1:0] matrixC9_5;
output [`DWIDTH-1:0] matrixC9_6;
output [`DWIDTH-1:0] matrixC9_7;
output [`DWIDTH-1:0] matrixC9_8;
output [`DWIDTH-1:0] matrixC9_9;
output [`DWIDTH-1:0] matrixC9_10;
output [`DWIDTH-1:0] matrixC9_11;
output [`DWIDTH-1:0] matrixC9_12;
output [`DWIDTH-1:0] matrixC9_13;
output [`DWIDTH-1:0] matrixC9_14;
output [`DWIDTH-1:0] matrixC9_15;
output [`DWIDTH-1:0] matrixC9_16;
output [`DWIDTH-1:0] matrixC9_17;
output [`DWIDTH-1:0] matrixC9_18;
output [`DWIDTH-1:0] matrixC9_19;
output [`DWIDTH-1:0] matrixC9_20;
output [`DWIDTH-1:0] matrixC9_21;
output [`DWIDTH-1:0] matrixC9_22;
output [`DWIDTH-1:0] matrixC9_23;
output [`DWIDTH-1:0] matrixC9_24;
output [`DWIDTH-1:0] matrixC9_25;
output [`DWIDTH-1:0] matrixC9_26;
output [`DWIDTH-1:0] matrixC9_27;
output [`DWIDTH-1:0] matrixC9_28;
output [`DWIDTH-1:0] matrixC9_29;
output [`DWIDTH-1:0] matrixC9_30;
output [`DWIDTH-1:0] matrixC9_31;
output [`DWIDTH-1:0] matrixC10_0;
output [`DWIDTH-1:0] matrixC10_1;
output [`DWIDTH-1:0] matrixC10_2;
output [`DWIDTH-1:0] matrixC10_3;
output [`DWIDTH-1:0] matrixC10_4;
output [`DWIDTH-1:0] matrixC10_5;
output [`DWIDTH-1:0] matrixC10_6;
output [`DWIDTH-1:0] matrixC10_7;
output [`DWIDTH-1:0] matrixC10_8;
output [`DWIDTH-1:0] matrixC10_9;
output [`DWIDTH-1:0] matrixC10_10;
output [`DWIDTH-1:0] matrixC10_11;
output [`DWIDTH-1:0] matrixC10_12;
output [`DWIDTH-1:0] matrixC10_13;
output [`DWIDTH-1:0] matrixC10_14;
output [`DWIDTH-1:0] matrixC10_15;
output [`DWIDTH-1:0] matrixC10_16;
output [`DWIDTH-1:0] matrixC10_17;
output [`DWIDTH-1:0] matrixC10_18;
output [`DWIDTH-1:0] matrixC10_19;
output [`DWIDTH-1:0] matrixC10_20;
output [`DWIDTH-1:0] matrixC10_21;
output [`DWIDTH-1:0] matrixC10_22;
output [`DWIDTH-1:0] matrixC10_23;
output [`DWIDTH-1:0] matrixC10_24;
output [`DWIDTH-1:0] matrixC10_25;
output [`DWIDTH-1:0] matrixC10_26;
output [`DWIDTH-1:0] matrixC10_27;
output [`DWIDTH-1:0] matrixC10_28;
output [`DWIDTH-1:0] matrixC10_29;
output [`DWIDTH-1:0] matrixC10_30;
output [`DWIDTH-1:0] matrixC10_31;
output [`DWIDTH-1:0] matrixC11_0;
output [`DWIDTH-1:0] matrixC11_1;
output [`DWIDTH-1:0] matrixC11_2;
output [`DWIDTH-1:0] matrixC11_3;
output [`DWIDTH-1:0] matrixC11_4;
output [`DWIDTH-1:0] matrixC11_5;
output [`DWIDTH-1:0] matrixC11_6;
output [`DWIDTH-1:0] matrixC11_7;
output [`DWIDTH-1:0] matrixC11_8;
output [`DWIDTH-1:0] matrixC11_9;
output [`DWIDTH-1:0] matrixC11_10;
output [`DWIDTH-1:0] matrixC11_11;
output [`DWIDTH-1:0] matrixC11_12;
output [`DWIDTH-1:0] matrixC11_13;
output [`DWIDTH-1:0] matrixC11_14;
output [`DWIDTH-1:0] matrixC11_15;
output [`DWIDTH-1:0] matrixC11_16;
output [`DWIDTH-1:0] matrixC11_17;
output [`DWIDTH-1:0] matrixC11_18;
output [`DWIDTH-1:0] matrixC11_19;
output [`DWIDTH-1:0] matrixC11_20;
output [`DWIDTH-1:0] matrixC11_21;
output [`DWIDTH-1:0] matrixC11_22;
output [`DWIDTH-1:0] matrixC11_23;
output [`DWIDTH-1:0] matrixC11_24;
output [`DWIDTH-1:0] matrixC11_25;
output [`DWIDTH-1:0] matrixC11_26;
output [`DWIDTH-1:0] matrixC11_27;
output [`DWIDTH-1:0] matrixC11_28;
output [`DWIDTH-1:0] matrixC11_29;
output [`DWIDTH-1:0] matrixC11_30;
output [`DWIDTH-1:0] matrixC11_31;
output [`DWIDTH-1:0] matrixC12_0;
output [`DWIDTH-1:0] matrixC12_1;
output [`DWIDTH-1:0] matrixC12_2;
output [`DWIDTH-1:0] matrixC12_3;
output [`DWIDTH-1:0] matrixC12_4;
output [`DWIDTH-1:0] matrixC12_5;
output [`DWIDTH-1:0] matrixC12_6;
output [`DWIDTH-1:0] matrixC12_7;
output [`DWIDTH-1:0] matrixC12_8;
output [`DWIDTH-1:0] matrixC12_9;
output [`DWIDTH-1:0] matrixC12_10;
output [`DWIDTH-1:0] matrixC12_11;
output [`DWIDTH-1:0] matrixC12_12;
output [`DWIDTH-1:0] matrixC12_13;
output [`DWIDTH-1:0] matrixC12_14;
output [`DWIDTH-1:0] matrixC12_15;
output [`DWIDTH-1:0] matrixC12_16;
output [`DWIDTH-1:0] matrixC12_17;
output [`DWIDTH-1:0] matrixC12_18;
output [`DWIDTH-1:0] matrixC12_19;
output [`DWIDTH-1:0] matrixC12_20;
output [`DWIDTH-1:0] matrixC12_21;
output [`DWIDTH-1:0] matrixC12_22;
output [`DWIDTH-1:0] matrixC12_23;
output [`DWIDTH-1:0] matrixC12_24;
output [`DWIDTH-1:0] matrixC12_25;
output [`DWIDTH-1:0] matrixC12_26;
output [`DWIDTH-1:0] matrixC12_27;
output [`DWIDTH-1:0] matrixC12_28;
output [`DWIDTH-1:0] matrixC12_29;
output [`DWIDTH-1:0] matrixC12_30;
output [`DWIDTH-1:0] matrixC12_31;
output [`DWIDTH-1:0] matrixC13_0;
output [`DWIDTH-1:0] matrixC13_1;
output [`DWIDTH-1:0] matrixC13_2;
output [`DWIDTH-1:0] matrixC13_3;
output [`DWIDTH-1:0] matrixC13_4;
output [`DWIDTH-1:0] matrixC13_5;
output [`DWIDTH-1:0] matrixC13_6;
output [`DWIDTH-1:0] matrixC13_7;
output [`DWIDTH-1:0] matrixC13_8;
output [`DWIDTH-1:0] matrixC13_9;
output [`DWIDTH-1:0] matrixC13_10;
output [`DWIDTH-1:0] matrixC13_11;
output [`DWIDTH-1:0] matrixC13_12;
output [`DWIDTH-1:0] matrixC13_13;
output [`DWIDTH-1:0] matrixC13_14;
output [`DWIDTH-1:0] matrixC13_15;
output [`DWIDTH-1:0] matrixC13_16;
output [`DWIDTH-1:0] matrixC13_17;
output [`DWIDTH-1:0] matrixC13_18;
output [`DWIDTH-1:0] matrixC13_19;
output [`DWIDTH-1:0] matrixC13_20;
output [`DWIDTH-1:0] matrixC13_21;
output [`DWIDTH-1:0] matrixC13_22;
output [`DWIDTH-1:0] matrixC13_23;
output [`DWIDTH-1:0] matrixC13_24;
output [`DWIDTH-1:0] matrixC13_25;
output [`DWIDTH-1:0] matrixC13_26;
output [`DWIDTH-1:0] matrixC13_27;
output [`DWIDTH-1:0] matrixC13_28;
output [`DWIDTH-1:0] matrixC13_29;
output [`DWIDTH-1:0] matrixC13_30;
output [`DWIDTH-1:0] matrixC13_31;
output [`DWIDTH-1:0] matrixC14_0;
output [`DWIDTH-1:0] matrixC14_1;
output [`DWIDTH-1:0] matrixC14_2;
output [`DWIDTH-1:0] matrixC14_3;
output [`DWIDTH-1:0] matrixC14_4;
output [`DWIDTH-1:0] matrixC14_5;
output [`DWIDTH-1:0] matrixC14_6;
output [`DWIDTH-1:0] matrixC14_7;
output [`DWIDTH-1:0] matrixC14_8;
output [`DWIDTH-1:0] matrixC14_9;
output [`DWIDTH-1:0] matrixC14_10;
output [`DWIDTH-1:0] matrixC14_11;
output [`DWIDTH-1:0] matrixC14_12;
output [`DWIDTH-1:0] matrixC14_13;
output [`DWIDTH-1:0] matrixC14_14;
output [`DWIDTH-1:0] matrixC14_15;
output [`DWIDTH-1:0] matrixC14_16;
output [`DWIDTH-1:0] matrixC14_17;
output [`DWIDTH-1:0] matrixC14_18;
output [`DWIDTH-1:0] matrixC14_19;
output [`DWIDTH-1:0] matrixC14_20;
output [`DWIDTH-1:0] matrixC14_21;
output [`DWIDTH-1:0] matrixC14_22;
output [`DWIDTH-1:0] matrixC14_23;
output [`DWIDTH-1:0] matrixC14_24;
output [`DWIDTH-1:0] matrixC14_25;
output [`DWIDTH-1:0] matrixC14_26;
output [`DWIDTH-1:0] matrixC14_27;
output [`DWIDTH-1:0] matrixC14_28;
output [`DWIDTH-1:0] matrixC14_29;
output [`DWIDTH-1:0] matrixC14_30;
output [`DWIDTH-1:0] matrixC14_31;
output [`DWIDTH-1:0] matrixC15_0;
output [`DWIDTH-1:0] matrixC15_1;
output [`DWIDTH-1:0] matrixC15_2;
output [`DWIDTH-1:0] matrixC15_3;
output [`DWIDTH-1:0] matrixC15_4;
output [`DWIDTH-1:0] matrixC15_5;
output [`DWIDTH-1:0] matrixC15_6;
output [`DWIDTH-1:0] matrixC15_7;
output [`DWIDTH-1:0] matrixC15_8;
output [`DWIDTH-1:0] matrixC15_9;
output [`DWIDTH-1:0] matrixC15_10;
output [`DWIDTH-1:0] matrixC15_11;
output [`DWIDTH-1:0] matrixC15_12;
output [`DWIDTH-1:0] matrixC15_13;
output [`DWIDTH-1:0] matrixC15_14;
output [`DWIDTH-1:0] matrixC15_15;
output [`DWIDTH-1:0] matrixC15_16;
output [`DWIDTH-1:0] matrixC15_17;
output [`DWIDTH-1:0] matrixC15_18;
output [`DWIDTH-1:0] matrixC15_19;
output [`DWIDTH-1:0] matrixC15_20;
output [`DWIDTH-1:0] matrixC15_21;
output [`DWIDTH-1:0] matrixC15_22;
output [`DWIDTH-1:0] matrixC15_23;
output [`DWIDTH-1:0] matrixC15_24;
output [`DWIDTH-1:0] matrixC15_25;
output [`DWIDTH-1:0] matrixC15_26;
output [`DWIDTH-1:0] matrixC15_27;
output [`DWIDTH-1:0] matrixC15_28;
output [`DWIDTH-1:0] matrixC15_29;
output [`DWIDTH-1:0] matrixC15_30;
output [`DWIDTH-1:0] matrixC15_31;
output [`DWIDTH-1:0] matrixC16_0;
output [`DWIDTH-1:0] matrixC16_1;
output [`DWIDTH-1:0] matrixC16_2;
output [`DWIDTH-1:0] matrixC16_3;
output [`DWIDTH-1:0] matrixC16_4;
output [`DWIDTH-1:0] matrixC16_5;
output [`DWIDTH-1:0] matrixC16_6;
output [`DWIDTH-1:0] matrixC16_7;
output [`DWIDTH-1:0] matrixC16_8;
output [`DWIDTH-1:0] matrixC16_9;
output [`DWIDTH-1:0] matrixC16_10;
output [`DWIDTH-1:0] matrixC16_11;
output [`DWIDTH-1:0] matrixC16_12;
output [`DWIDTH-1:0] matrixC16_13;
output [`DWIDTH-1:0] matrixC16_14;
output [`DWIDTH-1:0] matrixC16_15;
output [`DWIDTH-1:0] matrixC16_16;
output [`DWIDTH-1:0] matrixC16_17;
output [`DWIDTH-1:0] matrixC16_18;
output [`DWIDTH-1:0] matrixC16_19;
output [`DWIDTH-1:0] matrixC16_20;
output [`DWIDTH-1:0] matrixC16_21;
output [`DWIDTH-1:0] matrixC16_22;
output [`DWIDTH-1:0] matrixC16_23;
output [`DWIDTH-1:0] matrixC16_24;
output [`DWIDTH-1:0] matrixC16_25;
output [`DWIDTH-1:0] matrixC16_26;
output [`DWIDTH-1:0] matrixC16_27;
output [`DWIDTH-1:0] matrixC16_28;
output [`DWIDTH-1:0] matrixC16_29;
output [`DWIDTH-1:0] matrixC16_30;
output [`DWIDTH-1:0] matrixC16_31;
output [`DWIDTH-1:0] matrixC17_0;
output [`DWIDTH-1:0] matrixC17_1;
output [`DWIDTH-1:0] matrixC17_2;
output [`DWIDTH-1:0] matrixC17_3;
output [`DWIDTH-1:0] matrixC17_4;
output [`DWIDTH-1:0] matrixC17_5;
output [`DWIDTH-1:0] matrixC17_6;
output [`DWIDTH-1:0] matrixC17_7;
output [`DWIDTH-1:0] matrixC17_8;
output [`DWIDTH-1:0] matrixC17_9;
output [`DWIDTH-1:0] matrixC17_10;
output [`DWIDTH-1:0] matrixC17_11;
output [`DWIDTH-1:0] matrixC17_12;
output [`DWIDTH-1:0] matrixC17_13;
output [`DWIDTH-1:0] matrixC17_14;
output [`DWIDTH-1:0] matrixC17_15;
output [`DWIDTH-1:0] matrixC17_16;
output [`DWIDTH-1:0] matrixC17_17;
output [`DWIDTH-1:0] matrixC17_18;
output [`DWIDTH-1:0] matrixC17_19;
output [`DWIDTH-1:0] matrixC17_20;
output [`DWIDTH-1:0] matrixC17_21;
output [`DWIDTH-1:0] matrixC17_22;
output [`DWIDTH-1:0] matrixC17_23;
output [`DWIDTH-1:0] matrixC17_24;
output [`DWIDTH-1:0] matrixC17_25;
output [`DWIDTH-1:0] matrixC17_26;
output [`DWIDTH-1:0] matrixC17_27;
output [`DWIDTH-1:0] matrixC17_28;
output [`DWIDTH-1:0] matrixC17_29;
output [`DWIDTH-1:0] matrixC17_30;
output [`DWIDTH-1:0] matrixC17_31;
output [`DWIDTH-1:0] matrixC18_0;
output [`DWIDTH-1:0] matrixC18_1;
output [`DWIDTH-1:0] matrixC18_2;
output [`DWIDTH-1:0] matrixC18_3;
output [`DWIDTH-1:0] matrixC18_4;
output [`DWIDTH-1:0] matrixC18_5;
output [`DWIDTH-1:0] matrixC18_6;
output [`DWIDTH-1:0] matrixC18_7;
output [`DWIDTH-1:0] matrixC18_8;
output [`DWIDTH-1:0] matrixC18_9;
output [`DWIDTH-1:0] matrixC18_10;
output [`DWIDTH-1:0] matrixC18_11;
output [`DWIDTH-1:0] matrixC18_12;
output [`DWIDTH-1:0] matrixC18_13;
output [`DWIDTH-1:0] matrixC18_14;
output [`DWIDTH-1:0] matrixC18_15;
output [`DWIDTH-1:0] matrixC18_16;
output [`DWIDTH-1:0] matrixC18_17;
output [`DWIDTH-1:0] matrixC18_18;
output [`DWIDTH-1:0] matrixC18_19;
output [`DWIDTH-1:0] matrixC18_20;
output [`DWIDTH-1:0] matrixC18_21;
output [`DWIDTH-1:0] matrixC18_22;
output [`DWIDTH-1:0] matrixC18_23;
output [`DWIDTH-1:0] matrixC18_24;
output [`DWIDTH-1:0] matrixC18_25;
output [`DWIDTH-1:0] matrixC18_26;
output [`DWIDTH-1:0] matrixC18_27;
output [`DWIDTH-1:0] matrixC18_28;
output [`DWIDTH-1:0] matrixC18_29;
output [`DWIDTH-1:0] matrixC18_30;
output [`DWIDTH-1:0] matrixC18_31;
output [`DWIDTH-1:0] matrixC19_0;
output [`DWIDTH-1:0] matrixC19_1;
output [`DWIDTH-1:0] matrixC19_2;
output [`DWIDTH-1:0] matrixC19_3;
output [`DWIDTH-1:0] matrixC19_4;
output [`DWIDTH-1:0] matrixC19_5;
output [`DWIDTH-1:0] matrixC19_6;
output [`DWIDTH-1:0] matrixC19_7;
output [`DWIDTH-1:0] matrixC19_8;
output [`DWIDTH-1:0] matrixC19_9;
output [`DWIDTH-1:0] matrixC19_10;
output [`DWIDTH-1:0] matrixC19_11;
output [`DWIDTH-1:0] matrixC19_12;
output [`DWIDTH-1:0] matrixC19_13;
output [`DWIDTH-1:0] matrixC19_14;
output [`DWIDTH-1:0] matrixC19_15;
output [`DWIDTH-1:0] matrixC19_16;
output [`DWIDTH-1:0] matrixC19_17;
output [`DWIDTH-1:0] matrixC19_18;
output [`DWIDTH-1:0] matrixC19_19;
output [`DWIDTH-1:0] matrixC19_20;
output [`DWIDTH-1:0] matrixC19_21;
output [`DWIDTH-1:0] matrixC19_22;
output [`DWIDTH-1:0] matrixC19_23;
output [`DWIDTH-1:0] matrixC19_24;
output [`DWIDTH-1:0] matrixC19_25;
output [`DWIDTH-1:0] matrixC19_26;
output [`DWIDTH-1:0] matrixC19_27;
output [`DWIDTH-1:0] matrixC19_28;
output [`DWIDTH-1:0] matrixC19_29;
output [`DWIDTH-1:0] matrixC19_30;
output [`DWIDTH-1:0] matrixC19_31;
output [`DWIDTH-1:0] matrixC20_0;
output [`DWIDTH-1:0] matrixC20_1;
output [`DWIDTH-1:0] matrixC20_2;
output [`DWIDTH-1:0] matrixC20_3;
output [`DWIDTH-1:0] matrixC20_4;
output [`DWIDTH-1:0] matrixC20_5;
output [`DWIDTH-1:0] matrixC20_6;
output [`DWIDTH-1:0] matrixC20_7;
output [`DWIDTH-1:0] matrixC20_8;
output [`DWIDTH-1:0] matrixC20_9;
output [`DWIDTH-1:0] matrixC20_10;
output [`DWIDTH-1:0] matrixC20_11;
output [`DWIDTH-1:0] matrixC20_12;
output [`DWIDTH-1:0] matrixC20_13;
output [`DWIDTH-1:0] matrixC20_14;
output [`DWIDTH-1:0] matrixC20_15;
output [`DWIDTH-1:0] matrixC20_16;
output [`DWIDTH-1:0] matrixC20_17;
output [`DWIDTH-1:0] matrixC20_18;
output [`DWIDTH-1:0] matrixC20_19;
output [`DWIDTH-1:0] matrixC20_20;
output [`DWIDTH-1:0] matrixC20_21;
output [`DWIDTH-1:0] matrixC20_22;
output [`DWIDTH-1:0] matrixC20_23;
output [`DWIDTH-1:0] matrixC20_24;
output [`DWIDTH-1:0] matrixC20_25;
output [`DWIDTH-1:0] matrixC20_26;
output [`DWIDTH-1:0] matrixC20_27;
output [`DWIDTH-1:0] matrixC20_28;
output [`DWIDTH-1:0] matrixC20_29;
output [`DWIDTH-1:0] matrixC20_30;
output [`DWIDTH-1:0] matrixC20_31;
output [`DWIDTH-1:0] matrixC21_0;
output [`DWIDTH-1:0] matrixC21_1;
output [`DWIDTH-1:0] matrixC21_2;
output [`DWIDTH-1:0] matrixC21_3;
output [`DWIDTH-1:0] matrixC21_4;
output [`DWIDTH-1:0] matrixC21_5;
output [`DWIDTH-1:0] matrixC21_6;
output [`DWIDTH-1:0] matrixC21_7;
output [`DWIDTH-1:0] matrixC21_8;
output [`DWIDTH-1:0] matrixC21_9;
output [`DWIDTH-1:0] matrixC21_10;
output [`DWIDTH-1:0] matrixC21_11;
output [`DWIDTH-1:0] matrixC21_12;
output [`DWIDTH-1:0] matrixC21_13;
output [`DWIDTH-1:0] matrixC21_14;
output [`DWIDTH-1:0] matrixC21_15;
output [`DWIDTH-1:0] matrixC21_16;
output [`DWIDTH-1:0] matrixC21_17;
output [`DWIDTH-1:0] matrixC21_18;
output [`DWIDTH-1:0] matrixC21_19;
output [`DWIDTH-1:0] matrixC21_20;
output [`DWIDTH-1:0] matrixC21_21;
output [`DWIDTH-1:0] matrixC21_22;
output [`DWIDTH-1:0] matrixC21_23;
output [`DWIDTH-1:0] matrixC21_24;
output [`DWIDTH-1:0] matrixC21_25;
output [`DWIDTH-1:0] matrixC21_26;
output [`DWIDTH-1:0] matrixC21_27;
output [`DWIDTH-1:0] matrixC21_28;
output [`DWIDTH-1:0] matrixC21_29;
output [`DWIDTH-1:0] matrixC21_30;
output [`DWIDTH-1:0] matrixC21_31;
output [`DWIDTH-1:0] matrixC22_0;
output [`DWIDTH-1:0] matrixC22_1;
output [`DWIDTH-1:0] matrixC22_2;
output [`DWIDTH-1:0] matrixC22_3;
output [`DWIDTH-1:0] matrixC22_4;
output [`DWIDTH-1:0] matrixC22_5;
output [`DWIDTH-1:0] matrixC22_6;
output [`DWIDTH-1:0] matrixC22_7;
output [`DWIDTH-1:0] matrixC22_8;
output [`DWIDTH-1:0] matrixC22_9;
output [`DWIDTH-1:0] matrixC22_10;
output [`DWIDTH-1:0] matrixC22_11;
output [`DWIDTH-1:0] matrixC22_12;
output [`DWIDTH-1:0] matrixC22_13;
output [`DWIDTH-1:0] matrixC22_14;
output [`DWIDTH-1:0] matrixC22_15;
output [`DWIDTH-1:0] matrixC22_16;
output [`DWIDTH-1:0] matrixC22_17;
output [`DWIDTH-1:0] matrixC22_18;
output [`DWIDTH-1:0] matrixC22_19;
output [`DWIDTH-1:0] matrixC22_20;
output [`DWIDTH-1:0] matrixC22_21;
output [`DWIDTH-1:0] matrixC22_22;
output [`DWIDTH-1:0] matrixC22_23;
output [`DWIDTH-1:0] matrixC22_24;
output [`DWIDTH-1:0] matrixC22_25;
output [`DWIDTH-1:0] matrixC22_26;
output [`DWIDTH-1:0] matrixC22_27;
output [`DWIDTH-1:0] matrixC22_28;
output [`DWIDTH-1:0] matrixC22_29;
output [`DWIDTH-1:0] matrixC22_30;
output [`DWIDTH-1:0] matrixC22_31;
output [`DWIDTH-1:0] matrixC23_0;
output [`DWIDTH-1:0] matrixC23_1;
output [`DWIDTH-1:0] matrixC23_2;
output [`DWIDTH-1:0] matrixC23_3;
output [`DWIDTH-1:0] matrixC23_4;
output [`DWIDTH-1:0] matrixC23_5;
output [`DWIDTH-1:0] matrixC23_6;
output [`DWIDTH-1:0] matrixC23_7;
output [`DWIDTH-1:0] matrixC23_8;
output [`DWIDTH-1:0] matrixC23_9;
output [`DWIDTH-1:0] matrixC23_10;
output [`DWIDTH-1:0] matrixC23_11;
output [`DWIDTH-1:0] matrixC23_12;
output [`DWIDTH-1:0] matrixC23_13;
output [`DWIDTH-1:0] matrixC23_14;
output [`DWIDTH-1:0] matrixC23_15;
output [`DWIDTH-1:0] matrixC23_16;
output [`DWIDTH-1:0] matrixC23_17;
output [`DWIDTH-1:0] matrixC23_18;
output [`DWIDTH-1:0] matrixC23_19;
output [`DWIDTH-1:0] matrixC23_20;
output [`DWIDTH-1:0] matrixC23_21;
output [`DWIDTH-1:0] matrixC23_22;
output [`DWIDTH-1:0] matrixC23_23;
output [`DWIDTH-1:0] matrixC23_24;
output [`DWIDTH-1:0] matrixC23_25;
output [`DWIDTH-1:0] matrixC23_26;
output [`DWIDTH-1:0] matrixC23_27;
output [`DWIDTH-1:0] matrixC23_28;
output [`DWIDTH-1:0] matrixC23_29;
output [`DWIDTH-1:0] matrixC23_30;
output [`DWIDTH-1:0] matrixC23_31;
output [`DWIDTH-1:0] matrixC24_0;
output [`DWIDTH-1:0] matrixC24_1;
output [`DWIDTH-1:0] matrixC24_2;
output [`DWIDTH-1:0] matrixC24_3;
output [`DWIDTH-1:0] matrixC24_4;
output [`DWIDTH-1:0] matrixC24_5;
output [`DWIDTH-1:0] matrixC24_6;
output [`DWIDTH-1:0] matrixC24_7;
output [`DWIDTH-1:0] matrixC24_8;
output [`DWIDTH-1:0] matrixC24_9;
output [`DWIDTH-1:0] matrixC24_10;
output [`DWIDTH-1:0] matrixC24_11;
output [`DWIDTH-1:0] matrixC24_12;
output [`DWIDTH-1:0] matrixC24_13;
output [`DWIDTH-1:0] matrixC24_14;
output [`DWIDTH-1:0] matrixC24_15;
output [`DWIDTH-1:0] matrixC24_16;
output [`DWIDTH-1:0] matrixC24_17;
output [`DWIDTH-1:0] matrixC24_18;
output [`DWIDTH-1:0] matrixC24_19;
output [`DWIDTH-1:0] matrixC24_20;
output [`DWIDTH-1:0] matrixC24_21;
output [`DWIDTH-1:0] matrixC24_22;
output [`DWIDTH-1:0] matrixC24_23;
output [`DWIDTH-1:0] matrixC24_24;
output [`DWIDTH-1:0] matrixC24_25;
output [`DWIDTH-1:0] matrixC24_26;
output [`DWIDTH-1:0] matrixC24_27;
output [`DWIDTH-1:0] matrixC24_28;
output [`DWIDTH-1:0] matrixC24_29;
output [`DWIDTH-1:0] matrixC24_30;
output [`DWIDTH-1:0] matrixC24_31;
output [`DWIDTH-1:0] matrixC25_0;
output [`DWIDTH-1:0] matrixC25_1;
output [`DWIDTH-1:0] matrixC25_2;
output [`DWIDTH-1:0] matrixC25_3;
output [`DWIDTH-1:0] matrixC25_4;
output [`DWIDTH-1:0] matrixC25_5;
output [`DWIDTH-1:0] matrixC25_6;
output [`DWIDTH-1:0] matrixC25_7;
output [`DWIDTH-1:0] matrixC25_8;
output [`DWIDTH-1:0] matrixC25_9;
output [`DWIDTH-1:0] matrixC25_10;
output [`DWIDTH-1:0] matrixC25_11;
output [`DWIDTH-1:0] matrixC25_12;
output [`DWIDTH-1:0] matrixC25_13;
output [`DWIDTH-1:0] matrixC25_14;
output [`DWIDTH-1:0] matrixC25_15;
output [`DWIDTH-1:0] matrixC25_16;
output [`DWIDTH-1:0] matrixC25_17;
output [`DWIDTH-1:0] matrixC25_18;
output [`DWIDTH-1:0] matrixC25_19;
output [`DWIDTH-1:0] matrixC25_20;
output [`DWIDTH-1:0] matrixC25_21;
output [`DWIDTH-1:0] matrixC25_22;
output [`DWIDTH-1:0] matrixC25_23;
output [`DWIDTH-1:0] matrixC25_24;
output [`DWIDTH-1:0] matrixC25_25;
output [`DWIDTH-1:0] matrixC25_26;
output [`DWIDTH-1:0] matrixC25_27;
output [`DWIDTH-1:0] matrixC25_28;
output [`DWIDTH-1:0] matrixC25_29;
output [`DWIDTH-1:0] matrixC25_30;
output [`DWIDTH-1:0] matrixC25_31;
output [`DWIDTH-1:0] matrixC26_0;
output [`DWIDTH-1:0] matrixC26_1;
output [`DWIDTH-1:0] matrixC26_2;
output [`DWIDTH-1:0] matrixC26_3;
output [`DWIDTH-1:0] matrixC26_4;
output [`DWIDTH-1:0] matrixC26_5;
output [`DWIDTH-1:0] matrixC26_6;
output [`DWIDTH-1:0] matrixC26_7;
output [`DWIDTH-1:0] matrixC26_8;
output [`DWIDTH-1:0] matrixC26_9;
output [`DWIDTH-1:0] matrixC26_10;
output [`DWIDTH-1:0] matrixC26_11;
output [`DWIDTH-1:0] matrixC26_12;
output [`DWIDTH-1:0] matrixC26_13;
output [`DWIDTH-1:0] matrixC26_14;
output [`DWIDTH-1:0] matrixC26_15;
output [`DWIDTH-1:0] matrixC26_16;
output [`DWIDTH-1:0] matrixC26_17;
output [`DWIDTH-1:0] matrixC26_18;
output [`DWIDTH-1:0] matrixC26_19;
output [`DWIDTH-1:0] matrixC26_20;
output [`DWIDTH-1:0] matrixC26_21;
output [`DWIDTH-1:0] matrixC26_22;
output [`DWIDTH-1:0] matrixC26_23;
output [`DWIDTH-1:0] matrixC26_24;
output [`DWIDTH-1:0] matrixC26_25;
output [`DWIDTH-1:0] matrixC26_26;
output [`DWIDTH-1:0] matrixC26_27;
output [`DWIDTH-1:0] matrixC26_28;
output [`DWIDTH-1:0] matrixC26_29;
output [`DWIDTH-1:0] matrixC26_30;
output [`DWIDTH-1:0] matrixC26_31;
output [`DWIDTH-1:0] matrixC27_0;
output [`DWIDTH-1:0] matrixC27_1;
output [`DWIDTH-1:0] matrixC27_2;
output [`DWIDTH-1:0] matrixC27_3;
output [`DWIDTH-1:0] matrixC27_4;
output [`DWIDTH-1:0] matrixC27_5;
output [`DWIDTH-1:0] matrixC27_6;
output [`DWIDTH-1:0] matrixC27_7;
output [`DWIDTH-1:0] matrixC27_8;
output [`DWIDTH-1:0] matrixC27_9;
output [`DWIDTH-1:0] matrixC27_10;
output [`DWIDTH-1:0] matrixC27_11;
output [`DWIDTH-1:0] matrixC27_12;
output [`DWIDTH-1:0] matrixC27_13;
output [`DWIDTH-1:0] matrixC27_14;
output [`DWIDTH-1:0] matrixC27_15;
output [`DWIDTH-1:0] matrixC27_16;
output [`DWIDTH-1:0] matrixC27_17;
output [`DWIDTH-1:0] matrixC27_18;
output [`DWIDTH-1:0] matrixC27_19;
output [`DWIDTH-1:0] matrixC27_20;
output [`DWIDTH-1:0] matrixC27_21;
output [`DWIDTH-1:0] matrixC27_22;
output [`DWIDTH-1:0] matrixC27_23;
output [`DWIDTH-1:0] matrixC27_24;
output [`DWIDTH-1:0] matrixC27_25;
output [`DWIDTH-1:0] matrixC27_26;
output [`DWIDTH-1:0] matrixC27_27;
output [`DWIDTH-1:0] matrixC27_28;
output [`DWIDTH-1:0] matrixC27_29;
output [`DWIDTH-1:0] matrixC27_30;
output [`DWIDTH-1:0] matrixC27_31;
output [`DWIDTH-1:0] matrixC28_0;
output [`DWIDTH-1:0] matrixC28_1;
output [`DWIDTH-1:0] matrixC28_2;
output [`DWIDTH-1:0] matrixC28_3;
output [`DWIDTH-1:0] matrixC28_4;
output [`DWIDTH-1:0] matrixC28_5;
output [`DWIDTH-1:0] matrixC28_6;
output [`DWIDTH-1:0] matrixC28_7;
output [`DWIDTH-1:0] matrixC28_8;
output [`DWIDTH-1:0] matrixC28_9;
output [`DWIDTH-1:0] matrixC28_10;
output [`DWIDTH-1:0] matrixC28_11;
output [`DWIDTH-1:0] matrixC28_12;
output [`DWIDTH-1:0] matrixC28_13;
output [`DWIDTH-1:0] matrixC28_14;
output [`DWIDTH-1:0] matrixC28_15;
output [`DWIDTH-1:0] matrixC28_16;
output [`DWIDTH-1:0] matrixC28_17;
output [`DWIDTH-1:0] matrixC28_18;
output [`DWIDTH-1:0] matrixC28_19;
output [`DWIDTH-1:0] matrixC28_20;
output [`DWIDTH-1:0] matrixC28_21;
output [`DWIDTH-1:0] matrixC28_22;
output [`DWIDTH-1:0] matrixC28_23;
output [`DWIDTH-1:0] matrixC28_24;
output [`DWIDTH-1:0] matrixC28_25;
output [`DWIDTH-1:0] matrixC28_26;
output [`DWIDTH-1:0] matrixC28_27;
output [`DWIDTH-1:0] matrixC28_28;
output [`DWIDTH-1:0] matrixC28_29;
output [`DWIDTH-1:0] matrixC28_30;
output [`DWIDTH-1:0] matrixC28_31;
output [`DWIDTH-1:0] matrixC29_0;
output [`DWIDTH-1:0] matrixC29_1;
output [`DWIDTH-1:0] matrixC29_2;
output [`DWIDTH-1:0] matrixC29_3;
output [`DWIDTH-1:0] matrixC29_4;
output [`DWIDTH-1:0] matrixC29_5;
output [`DWIDTH-1:0] matrixC29_6;
output [`DWIDTH-1:0] matrixC29_7;
output [`DWIDTH-1:0] matrixC29_8;
output [`DWIDTH-1:0] matrixC29_9;
output [`DWIDTH-1:0] matrixC29_10;
output [`DWIDTH-1:0] matrixC29_11;
output [`DWIDTH-1:0] matrixC29_12;
output [`DWIDTH-1:0] matrixC29_13;
output [`DWIDTH-1:0] matrixC29_14;
output [`DWIDTH-1:0] matrixC29_15;
output [`DWIDTH-1:0] matrixC29_16;
output [`DWIDTH-1:0] matrixC29_17;
output [`DWIDTH-1:0] matrixC29_18;
output [`DWIDTH-1:0] matrixC29_19;
output [`DWIDTH-1:0] matrixC29_20;
output [`DWIDTH-1:0] matrixC29_21;
output [`DWIDTH-1:0] matrixC29_22;
output [`DWIDTH-1:0] matrixC29_23;
output [`DWIDTH-1:0] matrixC29_24;
output [`DWIDTH-1:0] matrixC29_25;
output [`DWIDTH-1:0] matrixC29_26;
output [`DWIDTH-1:0] matrixC29_27;
output [`DWIDTH-1:0] matrixC29_28;
output [`DWIDTH-1:0] matrixC29_29;
output [`DWIDTH-1:0] matrixC29_30;
output [`DWIDTH-1:0] matrixC29_31;
output [`DWIDTH-1:0] matrixC30_0;
output [`DWIDTH-1:0] matrixC30_1;
output [`DWIDTH-1:0] matrixC30_2;
output [`DWIDTH-1:0] matrixC30_3;
output [`DWIDTH-1:0] matrixC30_4;
output [`DWIDTH-1:0] matrixC30_5;
output [`DWIDTH-1:0] matrixC30_6;
output [`DWIDTH-1:0] matrixC30_7;
output [`DWIDTH-1:0] matrixC30_8;
output [`DWIDTH-1:0] matrixC30_9;
output [`DWIDTH-1:0] matrixC30_10;
output [`DWIDTH-1:0] matrixC30_11;
output [`DWIDTH-1:0] matrixC30_12;
output [`DWIDTH-1:0] matrixC30_13;
output [`DWIDTH-1:0] matrixC30_14;
output [`DWIDTH-1:0] matrixC30_15;
output [`DWIDTH-1:0] matrixC30_16;
output [`DWIDTH-1:0] matrixC30_17;
output [`DWIDTH-1:0] matrixC30_18;
output [`DWIDTH-1:0] matrixC30_19;
output [`DWIDTH-1:0] matrixC30_20;
output [`DWIDTH-1:0] matrixC30_21;
output [`DWIDTH-1:0] matrixC30_22;
output [`DWIDTH-1:0] matrixC30_23;
output [`DWIDTH-1:0] matrixC30_24;
output [`DWIDTH-1:0] matrixC30_25;
output [`DWIDTH-1:0] matrixC30_26;
output [`DWIDTH-1:0] matrixC30_27;
output [`DWIDTH-1:0] matrixC30_28;
output [`DWIDTH-1:0] matrixC30_29;
output [`DWIDTH-1:0] matrixC30_30;
output [`DWIDTH-1:0] matrixC30_31;
output [`DWIDTH-1:0] matrixC31_0;
output [`DWIDTH-1:0] matrixC31_1;
output [`DWIDTH-1:0] matrixC31_2;
output [`DWIDTH-1:0] matrixC31_3;
output [`DWIDTH-1:0] matrixC31_4;
output [`DWIDTH-1:0] matrixC31_5;
output [`DWIDTH-1:0] matrixC31_6;
output [`DWIDTH-1:0] matrixC31_7;
output [`DWIDTH-1:0] matrixC31_8;
output [`DWIDTH-1:0] matrixC31_9;
output [`DWIDTH-1:0] matrixC31_10;
output [`DWIDTH-1:0] matrixC31_11;
output [`DWIDTH-1:0] matrixC31_12;
output [`DWIDTH-1:0] matrixC31_13;
output [`DWIDTH-1:0] matrixC31_14;
output [`DWIDTH-1:0] matrixC31_15;
output [`DWIDTH-1:0] matrixC31_16;
output [`DWIDTH-1:0] matrixC31_17;
output [`DWIDTH-1:0] matrixC31_18;
output [`DWIDTH-1:0] matrixC31_19;
output [`DWIDTH-1:0] matrixC31_20;
output [`DWIDTH-1:0] matrixC31_21;
output [`DWIDTH-1:0] matrixC31_22;
output [`DWIDTH-1:0] matrixC31_23;
output [`DWIDTH-1:0] matrixC31_24;
output [`DWIDTH-1:0] matrixC31_25;
output [`DWIDTH-1:0] matrixC31_26;
output [`DWIDTH-1:0] matrixC31_27;
output [`DWIDTH-1:0] matrixC31_28;
output [`DWIDTH-1:0] matrixC31_29;
output [`DWIDTH-1:0] matrixC31_30;
output [`DWIDTH-1:0] matrixC31_31;

output [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data_out;
output [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data_out;

wire [`DWIDTH-1:0] a0_0to0_1, a0_1to0_2, a0_2to0_3, a0_3to0_4, a0_4to0_5, a0_5to0_6, a0_6to0_7, a0_7to0_8, a0_8to0_9, a0_9to0_10, a0_10to0_11, a0_11to0_12, a0_12to0_13, a0_13to0_14, a0_14to0_15, a0_15to0_16, a0_16to0_17, a0_17to0_18, a0_18to0_19, a0_19to0_20, a0_20to0_21, a0_21to0_22, a0_22to0_23, a0_23to0_24, a0_24to0_25, a0_25to0_26, a0_26to0_27, a0_27to0_28, a0_28to0_29, a0_29to0_30, a0_30to0_31, a0_31to0_32;
wire [`DWIDTH-1:0] a1_0to1_1, a1_1to1_2, a1_2to1_3, a1_3to1_4, a1_4to1_5, a1_5to1_6, a1_6to1_7, a1_7to1_8, a1_8to1_9, a1_9to1_10, a1_10to1_11, a1_11to1_12, a1_12to1_13, a1_13to1_14, a1_14to1_15, a1_15to1_16, a1_16to1_17, a1_17to1_18, a1_18to1_19, a1_19to1_20, a1_20to1_21, a1_21to1_22, a1_22to1_23, a1_23to1_24, a1_24to1_25, a1_25to1_26, a1_26to1_27, a1_27to1_28, a1_28to1_29, a1_29to1_30, a1_30to1_31, a1_31to1_32;
wire [`DWIDTH-1:0] a2_0to2_1, a2_1to2_2, a2_2to2_3, a2_3to2_4, a2_4to2_5, a2_5to2_6, a2_6to2_7, a2_7to2_8, a2_8to2_9, a2_9to2_10, a2_10to2_11, a2_11to2_12, a2_12to2_13, a2_13to2_14, a2_14to2_15, a2_15to2_16, a2_16to2_17, a2_17to2_18, a2_18to2_19, a2_19to2_20, a2_20to2_21, a2_21to2_22, a2_22to2_23, a2_23to2_24, a2_24to2_25, a2_25to2_26, a2_26to2_27, a2_27to2_28, a2_28to2_29, a2_29to2_30, a2_30to2_31, a2_31to2_32;
wire [`DWIDTH-1:0] a3_0to3_1, a3_1to3_2, a3_2to3_3, a3_3to3_4, a3_4to3_5, a3_5to3_6, a3_6to3_7, a3_7to3_8, a3_8to3_9, a3_9to3_10, a3_10to3_11, a3_11to3_12, a3_12to3_13, a3_13to3_14, a3_14to3_15, a3_15to3_16, a3_16to3_17, a3_17to3_18, a3_18to3_19, a3_19to3_20, a3_20to3_21, a3_21to3_22, a3_22to3_23, a3_23to3_24, a3_24to3_25, a3_25to3_26, a3_26to3_27, a3_27to3_28, a3_28to3_29, a3_29to3_30, a3_30to3_31, a3_31to3_32;
wire [`DWIDTH-1:0] a4_0to4_1, a4_1to4_2, a4_2to4_3, a4_3to4_4, a4_4to4_5, a4_5to4_6, a4_6to4_7, a4_7to4_8, a4_8to4_9, a4_9to4_10, a4_10to4_11, a4_11to4_12, a4_12to4_13, a4_13to4_14, a4_14to4_15, a4_15to4_16, a4_16to4_17, a4_17to4_18, a4_18to4_19, a4_19to4_20, a4_20to4_21, a4_21to4_22, a4_22to4_23, a4_23to4_24, a4_24to4_25, a4_25to4_26, a4_26to4_27, a4_27to4_28, a4_28to4_29, a4_29to4_30, a4_30to4_31, a4_31to4_32;
wire [`DWIDTH-1:0] a5_0to5_1, a5_1to5_2, a5_2to5_3, a5_3to5_4, a5_4to5_5, a5_5to5_6, a5_6to5_7, a5_7to5_8, a5_8to5_9, a5_9to5_10, a5_10to5_11, a5_11to5_12, a5_12to5_13, a5_13to5_14, a5_14to5_15, a5_15to5_16, a5_16to5_17, a5_17to5_18, a5_18to5_19, a5_19to5_20, a5_20to5_21, a5_21to5_22, a5_22to5_23, a5_23to5_24, a5_24to5_25, a5_25to5_26, a5_26to5_27, a5_27to5_28, a5_28to5_29, a5_29to5_30, a5_30to5_31, a5_31to5_32;
wire [`DWIDTH-1:0] a6_0to6_1, a6_1to6_2, a6_2to6_3, a6_3to6_4, a6_4to6_5, a6_5to6_6, a6_6to6_7, a6_7to6_8, a6_8to6_9, a6_9to6_10, a6_10to6_11, a6_11to6_12, a6_12to6_13, a6_13to6_14, a6_14to6_15, a6_15to6_16, a6_16to6_17, a6_17to6_18, a6_18to6_19, a6_19to6_20, a6_20to6_21, a6_21to6_22, a6_22to6_23, a6_23to6_24, a6_24to6_25, a6_25to6_26, a6_26to6_27, a6_27to6_28, a6_28to6_29, a6_29to6_30, a6_30to6_31, a6_31to6_32;
wire [`DWIDTH-1:0] a7_0to7_1, a7_1to7_2, a7_2to7_3, a7_3to7_4, a7_4to7_5, a7_5to7_6, a7_6to7_7, a7_7to7_8, a7_8to7_9, a7_9to7_10, a7_10to7_11, a7_11to7_12, a7_12to7_13, a7_13to7_14, a7_14to7_15, a7_15to7_16, a7_16to7_17, a7_17to7_18, a7_18to7_19, a7_19to7_20, a7_20to7_21, a7_21to7_22, a7_22to7_23, a7_23to7_24, a7_24to7_25, a7_25to7_26, a7_26to7_27, a7_27to7_28, a7_28to7_29, a7_29to7_30, a7_30to7_31, a7_31to7_32;
wire [`DWIDTH-1:0] a8_0to8_1, a8_1to8_2, a8_2to8_3, a8_3to8_4, a8_4to8_5, a8_5to8_6, a8_6to8_7, a8_7to8_8, a8_8to8_9, a8_9to8_10, a8_10to8_11, a8_11to8_12, a8_12to8_13, a8_13to8_14, a8_14to8_15, a8_15to8_16, a8_16to8_17, a8_17to8_18, a8_18to8_19, a8_19to8_20, a8_20to8_21, a8_21to8_22, a8_22to8_23, a8_23to8_24, a8_24to8_25, a8_25to8_26, a8_26to8_27, a8_27to8_28, a8_28to8_29, a8_29to8_30, a8_30to8_31, a8_31to8_32;
wire [`DWIDTH-1:0] a9_0to9_1, a9_1to9_2, a9_2to9_3, a9_3to9_4, a9_4to9_5, a9_5to9_6, a9_6to9_7, a9_7to9_8, a9_8to9_9, a9_9to9_10, a9_10to9_11, a9_11to9_12, a9_12to9_13, a9_13to9_14, a9_14to9_15, a9_15to9_16, a9_16to9_17, a9_17to9_18, a9_18to9_19, a9_19to9_20, a9_20to9_21, a9_21to9_22, a9_22to9_23, a9_23to9_24, a9_24to9_25, a9_25to9_26, a9_26to9_27, a9_27to9_28, a9_28to9_29, a9_29to9_30, a9_30to9_31, a9_31to9_32;
wire [`DWIDTH-1:0] a10_0to10_1, a10_1to10_2, a10_2to10_3, a10_3to10_4, a10_4to10_5, a10_5to10_6, a10_6to10_7, a10_7to10_8, a10_8to10_9, a10_9to10_10, a10_10to10_11, a10_11to10_12, a10_12to10_13, a10_13to10_14, a10_14to10_15, a10_15to10_16, a10_16to10_17, a10_17to10_18, a10_18to10_19, a10_19to10_20, a10_20to10_21, a10_21to10_22, a10_22to10_23, a10_23to10_24, a10_24to10_25, a10_25to10_26, a10_26to10_27, a10_27to10_28, a10_28to10_29, a10_29to10_30, a10_30to10_31, a10_31to10_32;
wire [`DWIDTH-1:0] a11_0to11_1, a11_1to11_2, a11_2to11_3, a11_3to11_4, a11_4to11_5, a11_5to11_6, a11_6to11_7, a11_7to11_8, a11_8to11_9, a11_9to11_10, a11_10to11_11, a11_11to11_12, a11_12to11_13, a11_13to11_14, a11_14to11_15, a11_15to11_16, a11_16to11_17, a11_17to11_18, a11_18to11_19, a11_19to11_20, a11_20to11_21, a11_21to11_22, a11_22to11_23, a11_23to11_24, a11_24to11_25, a11_25to11_26, a11_26to11_27, a11_27to11_28, a11_28to11_29, a11_29to11_30, a11_30to11_31, a11_31to11_32;
wire [`DWIDTH-1:0] a12_0to12_1, a12_1to12_2, a12_2to12_3, a12_3to12_4, a12_4to12_5, a12_5to12_6, a12_6to12_7, a12_7to12_8, a12_8to12_9, a12_9to12_10, a12_10to12_11, a12_11to12_12, a12_12to12_13, a12_13to12_14, a12_14to12_15, a12_15to12_16, a12_16to12_17, a12_17to12_18, a12_18to12_19, a12_19to12_20, a12_20to12_21, a12_21to12_22, a12_22to12_23, a12_23to12_24, a12_24to12_25, a12_25to12_26, a12_26to12_27, a12_27to12_28, a12_28to12_29, a12_29to12_30, a12_30to12_31, a12_31to12_32;
wire [`DWIDTH-1:0] a13_0to13_1, a13_1to13_2, a13_2to13_3, a13_3to13_4, a13_4to13_5, a13_5to13_6, a13_6to13_7, a13_7to13_8, a13_8to13_9, a13_9to13_10, a13_10to13_11, a13_11to13_12, a13_12to13_13, a13_13to13_14, a13_14to13_15, a13_15to13_16, a13_16to13_17, a13_17to13_18, a13_18to13_19, a13_19to13_20, a13_20to13_21, a13_21to13_22, a13_22to13_23, a13_23to13_24, a13_24to13_25, a13_25to13_26, a13_26to13_27, a13_27to13_28, a13_28to13_29, a13_29to13_30, a13_30to13_31, a13_31to13_32;
wire [`DWIDTH-1:0] a14_0to14_1, a14_1to14_2, a14_2to14_3, a14_3to14_4, a14_4to14_5, a14_5to14_6, a14_6to14_7, a14_7to14_8, a14_8to14_9, a14_9to14_10, a14_10to14_11, a14_11to14_12, a14_12to14_13, a14_13to14_14, a14_14to14_15, a14_15to14_16, a14_16to14_17, a14_17to14_18, a14_18to14_19, a14_19to14_20, a14_20to14_21, a14_21to14_22, a14_22to14_23, a14_23to14_24, a14_24to14_25, a14_25to14_26, a14_26to14_27, a14_27to14_28, a14_28to14_29, a14_29to14_30, a14_30to14_31, a14_31to14_32;
wire [`DWIDTH-1:0] a15_0to15_1, a15_1to15_2, a15_2to15_3, a15_3to15_4, a15_4to15_5, a15_5to15_6, a15_6to15_7, a15_7to15_8, a15_8to15_9, a15_9to15_10, a15_10to15_11, a15_11to15_12, a15_12to15_13, a15_13to15_14, a15_14to15_15, a15_15to15_16, a15_16to15_17, a15_17to15_18, a15_18to15_19, a15_19to15_20, a15_20to15_21, a15_21to15_22, a15_22to15_23, a15_23to15_24, a15_24to15_25, a15_25to15_26, a15_26to15_27, a15_27to15_28, a15_28to15_29, a15_29to15_30, a15_30to15_31, a15_31to15_32;
wire [`DWIDTH-1:0] a16_0to16_1, a16_1to16_2, a16_2to16_3, a16_3to16_4, a16_4to16_5, a16_5to16_6, a16_6to16_7, a16_7to16_8, a16_8to16_9, a16_9to16_10, a16_10to16_11, a16_11to16_12, a16_12to16_13, a16_13to16_14, a16_14to16_15, a16_15to16_16, a16_16to16_17, a16_17to16_18, a16_18to16_19, a16_19to16_20, a16_20to16_21, a16_21to16_22, a16_22to16_23, a16_23to16_24, a16_24to16_25, a16_25to16_26, a16_26to16_27, a16_27to16_28, a16_28to16_29, a16_29to16_30, a16_30to16_31, a16_31to16_32;
wire [`DWIDTH-1:0] a17_0to17_1, a17_1to17_2, a17_2to17_3, a17_3to17_4, a17_4to17_5, a17_5to17_6, a17_6to17_7, a17_7to17_8, a17_8to17_9, a17_9to17_10, a17_10to17_11, a17_11to17_12, a17_12to17_13, a17_13to17_14, a17_14to17_15, a17_15to17_16, a17_16to17_17, a17_17to17_18, a17_18to17_19, a17_19to17_20, a17_20to17_21, a17_21to17_22, a17_22to17_23, a17_23to17_24, a17_24to17_25, a17_25to17_26, a17_26to17_27, a17_27to17_28, a17_28to17_29, a17_29to17_30, a17_30to17_31, a17_31to17_32;
wire [`DWIDTH-1:0] a18_0to18_1, a18_1to18_2, a18_2to18_3, a18_3to18_4, a18_4to18_5, a18_5to18_6, a18_6to18_7, a18_7to18_8, a18_8to18_9, a18_9to18_10, a18_10to18_11, a18_11to18_12, a18_12to18_13, a18_13to18_14, a18_14to18_15, a18_15to18_16, a18_16to18_17, a18_17to18_18, a18_18to18_19, a18_19to18_20, a18_20to18_21, a18_21to18_22, a18_22to18_23, a18_23to18_24, a18_24to18_25, a18_25to18_26, a18_26to18_27, a18_27to18_28, a18_28to18_29, a18_29to18_30, a18_30to18_31, a18_31to18_32;
wire [`DWIDTH-1:0] a19_0to19_1, a19_1to19_2, a19_2to19_3, a19_3to19_4, a19_4to19_5, a19_5to19_6, a19_6to19_7, a19_7to19_8, a19_8to19_9, a19_9to19_10, a19_10to19_11, a19_11to19_12, a19_12to19_13, a19_13to19_14, a19_14to19_15, a19_15to19_16, a19_16to19_17, a19_17to19_18, a19_18to19_19, a19_19to19_20, a19_20to19_21, a19_21to19_22, a19_22to19_23, a19_23to19_24, a19_24to19_25, a19_25to19_26, a19_26to19_27, a19_27to19_28, a19_28to19_29, a19_29to19_30, a19_30to19_31, a19_31to19_32;
wire [`DWIDTH-1:0] a20_0to20_1, a20_1to20_2, a20_2to20_3, a20_3to20_4, a20_4to20_5, a20_5to20_6, a20_6to20_7, a20_7to20_8, a20_8to20_9, a20_9to20_10, a20_10to20_11, a20_11to20_12, a20_12to20_13, a20_13to20_14, a20_14to20_15, a20_15to20_16, a20_16to20_17, a20_17to20_18, a20_18to20_19, a20_19to20_20, a20_20to20_21, a20_21to20_22, a20_22to20_23, a20_23to20_24, a20_24to20_25, a20_25to20_26, a20_26to20_27, a20_27to20_28, a20_28to20_29, a20_29to20_30, a20_30to20_31, a20_31to20_32;
wire [`DWIDTH-1:0] a21_0to21_1, a21_1to21_2, a21_2to21_3, a21_3to21_4, a21_4to21_5, a21_5to21_6, a21_6to21_7, a21_7to21_8, a21_8to21_9, a21_9to21_10, a21_10to21_11, a21_11to21_12, a21_12to21_13, a21_13to21_14, a21_14to21_15, a21_15to21_16, a21_16to21_17, a21_17to21_18, a21_18to21_19, a21_19to21_20, a21_20to21_21, a21_21to21_22, a21_22to21_23, a21_23to21_24, a21_24to21_25, a21_25to21_26, a21_26to21_27, a21_27to21_28, a21_28to21_29, a21_29to21_30, a21_30to21_31, a21_31to21_32;
wire [`DWIDTH-1:0] a22_0to22_1, a22_1to22_2, a22_2to22_3, a22_3to22_4, a22_4to22_5, a22_5to22_6, a22_6to22_7, a22_7to22_8, a22_8to22_9, a22_9to22_10, a22_10to22_11, a22_11to22_12, a22_12to22_13, a22_13to22_14, a22_14to22_15, a22_15to22_16, a22_16to22_17, a22_17to22_18, a22_18to22_19, a22_19to22_20, a22_20to22_21, a22_21to22_22, a22_22to22_23, a22_23to22_24, a22_24to22_25, a22_25to22_26, a22_26to22_27, a22_27to22_28, a22_28to22_29, a22_29to22_30, a22_30to22_31, a22_31to22_32;
wire [`DWIDTH-1:0] a23_0to23_1, a23_1to23_2, a23_2to23_3, a23_3to23_4, a23_4to23_5, a23_5to23_6, a23_6to23_7, a23_7to23_8, a23_8to23_9, a23_9to23_10, a23_10to23_11, a23_11to23_12, a23_12to23_13, a23_13to23_14, a23_14to23_15, a23_15to23_16, a23_16to23_17, a23_17to23_18, a23_18to23_19, a23_19to23_20, a23_20to23_21, a23_21to23_22, a23_22to23_23, a23_23to23_24, a23_24to23_25, a23_25to23_26, a23_26to23_27, a23_27to23_28, a23_28to23_29, a23_29to23_30, a23_30to23_31, a23_31to23_32;
wire [`DWIDTH-1:0] a24_0to24_1, a24_1to24_2, a24_2to24_3, a24_3to24_4, a24_4to24_5, a24_5to24_6, a24_6to24_7, a24_7to24_8, a24_8to24_9, a24_9to24_10, a24_10to24_11, a24_11to24_12, a24_12to24_13, a24_13to24_14, a24_14to24_15, a24_15to24_16, a24_16to24_17, a24_17to24_18, a24_18to24_19, a24_19to24_20, a24_20to24_21, a24_21to24_22, a24_22to24_23, a24_23to24_24, a24_24to24_25, a24_25to24_26, a24_26to24_27, a24_27to24_28, a24_28to24_29, a24_29to24_30, a24_30to24_31, a24_31to24_32;
wire [`DWIDTH-1:0] a25_0to25_1, a25_1to25_2, a25_2to25_3, a25_3to25_4, a25_4to25_5, a25_5to25_6, a25_6to25_7, a25_7to25_8, a25_8to25_9, a25_9to25_10, a25_10to25_11, a25_11to25_12, a25_12to25_13, a25_13to25_14, a25_14to25_15, a25_15to25_16, a25_16to25_17, a25_17to25_18, a25_18to25_19, a25_19to25_20, a25_20to25_21, a25_21to25_22, a25_22to25_23, a25_23to25_24, a25_24to25_25, a25_25to25_26, a25_26to25_27, a25_27to25_28, a25_28to25_29, a25_29to25_30, a25_30to25_31, a25_31to25_32;
wire [`DWIDTH-1:0] a26_0to26_1, a26_1to26_2, a26_2to26_3, a26_3to26_4, a26_4to26_5, a26_5to26_6, a26_6to26_7, a26_7to26_8, a26_8to26_9, a26_9to26_10, a26_10to26_11, a26_11to26_12, a26_12to26_13, a26_13to26_14, a26_14to26_15, a26_15to26_16, a26_16to26_17, a26_17to26_18, a26_18to26_19, a26_19to26_20, a26_20to26_21, a26_21to26_22, a26_22to26_23, a26_23to26_24, a26_24to26_25, a26_25to26_26, a26_26to26_27, a26_27to26_28, a26_28to26_29, a26_29to26_30, a26_30to26_31, a26_31to26_32;
wire [`DWIDTH-1:0] a27_0to27_1, a27_1to27_2, a27_2to27_3, a27_3to27_4, a27_4to27_5, a27_5to27_6, a27_6to27_7, a27_7to27_8, a27_8to27_9, a27_9to27_10, a27_10to27_11, a27_11to27_12, a27_12to27_13, a27_13to27_14, a27_14to27_15, a27_15to27_16, a27_16to27_17, a27_17to27_18, a27_18to27_19, a27_19to27_20, a27_20to27_21, a27_21to27_22, a27_22to27_23, a27_23to27_24, a27_24to27_25, a27_25to27_26, a27_26to27_27, a27_27to27_28, a27_28to27_29, a27_29to27_30, a27_30to27_31, a27_31to27_32;
wire [`DWIDTH-1:0] a28_0to28_1, a28_1to28_2, a28_2to28_3, a28_3to28_4, a28_4to28_5, a28_5to28_6, a28_6to28_7, a28_7to28_8, a28_8to28_9, a28_9to28_10, a28_10to28_11, a28_11to28_12, a28_12to28_13, a28_13to28_14, a28_14to28_15, a28_15to28_16, a28_16to28_17, a28_17to28_18, a28_18to28_19, a28_19to28_20, a28_20to28_21, a28_21to28_22, a28_22to28_23, a28_23to28_24, a28_24to28_25, a28_25to28_26, a28_26to28_27, a28_27to28_28, a28_28to28_29, a28_29to28_30, a28_30to28_31, a28_31to28_32;
wire [`DWIDTH-1:0] a29_0to29_1, a29_1to29_2, a29_2to29_3, a29_3to29_4, a29_4to29_5, a29_5to29_6, a29_6to29_7, a29_7to29_8, a29_8to29_9, a29_9to29_10, a29_10to29_11, a29_11to29_12, a29_12to29_13, a29_13to29_14, a29_14to29_15, a29_15to29_16, a29_16to29_17, a29_17to29_18, a29_18to29_19, a29_19to29_20, a29_20to29_21, a29_21to29_22, a29_22to29_23, a29_23to29_24, a29_24to29_25, a29_25to29_26, a29_26to29_27, a29_27to29_28, a29_28to29_29, a29_29to29_30, a29_30to29_31, a29_31to29_32;
wire [`DWIDTH-1:0] a30_0to30_1, a30_1to30_2, a30_2to30_3, a30_3to30_4, a30_4to30_5, a30_5to30_6, a30_6to30_7, a30_7to30_8, a30_8to30_9, a30_9to30_10, a30_10to30_11, a30_11to30_12, a30_12to30_13, a30_13to30_14, a30_14to30_15, a30_15to30_16, a30_16to30_17, a30_17to30_18, a30_18to30_19, a30_19to30_20, a30_20to30_21, a30_21to30_22, a30_22to30_23, a30_23to30_24, a30_24to30_25, a30_25to30_26, a30_26to30_27, a30_27to30_28, a30_28to30_29, a30_29to30_30, a30_30to30_31, a30_31to30_32;
wire [`DWIDTH-1:0] a31_0to31_1, a31_1to31_2, a31_2to31_3, a31_3to31_4, a31_4to31_5, a31_5to31_6, a31_6to31_7, a31_7to31_8, a31_8to31_9, a31_9to31_10, a31_10to31_11, a31_11to31_12, a31_12to31_13, a31_13to31_14, a31_14to31_15, a31_15to31_16, a31_16to31_17, a31_17to31_18, a31_18to31_19, a31_19to31_20, a31_20to31_21, a31_21to31_22, a31_22to31_23, a31_23to31_24, a31_24to31_25, a31_25to31_26, a31_26to31_27, a31_27to31_28, a31_28to31_29, a31_29to31_30, a31_30to31_31, a31_31to31_32;

wire [`DWIDTH-1:0] b0_0to1_0, b1_0to2_0, b2_0to3_0, b3_0to4_0, b4_0to5_0, b5_0to6_0, b6_0to7_0, b7_0to8_0, b8_0to9_0, b9_0to10_0, b10_0to11_0, b11_0to12_0, b12_0to13_0, b13_0to14_0, b14_0to15_0, b15_0to16_0, b16_0to17_0, b17_0to18_0, b18_0to19_0, b19_0to20_0, b20_0to21_0, b21_0to22_0, b22_0to23_0, b23_0to24_0, b24_0to25_0, b25_0to26_0, b26_0to27_0, b27_0to28_0, b28_0to29_0, b29_0to30_0, b30_0to31_0, b31_0to32_0;
wire [`DWIDTH-1:0] b0_1to1_1, b1_1to2_1, b2_1to3_1, b3_1to4_1, b4_1to5_1, b5_1to6_1, b6_1to7_1, b7_1to8_1, b8_1to9_1, b9_1to10_1, b10_1to11_1, b11_1to12_1, b12_1to13_1, b13_1to14_1, b14_1to15_1, b15_1to16_1, b16_1to17_1, b17_1to18_1, b18_1to19_1, b19_1to20_1, b20_1to21_1, b21_1to22_1, b22_1to23_1, b23_1to24_1, b24_1to25_1, b25_1to26_1, b26_1to27_1, b27_1to28_1, b28_1to29_1, b29_1to30_1, b30_1to31_1, b31_1to32_1;
wire [`DWIDTH-1:0] b0_2to1_2, b1_2to2_2, b2_2to3_2, b3_2to4_2, b4_2to5_2, b5_2to6_2, b6_2to7_2, b7_2to8_2, b8_2to9_2, b9_2to10_2, b10_2to11_2, b11_2to12_2, b12_2to13_2, b13_2to14_2, b14_2to15_2, b15_2to16_2, b16_2to17_2, b17_2to18_2, b18_2to19_2, b19_2to20_2, b20_2to21_2, b21_2to22_2, b22_2to23_2, b23_2to24_2, b24_2to25_2, b25_2to26_2, b26_2to27_2, b27_2to28_2, b28_2to29_2, b29_2to30_2, b30_2to31_2, b31_2to32_2;
wire [`DWIDTH-1:0] b0_3to1_3, b1_3to2_3, b2_3to3_3, b3_3to4_3, b4_3to5_3, b5_3to6_3, b6_3to7_3, b7_3to8_3, b8_3to9_3, b9_3to10_3, b10_3to11_3, b11_3to12_3, b12_3to13_3, b13_3to14_3, b14_3to15_3, b15_3to16_3, b16_3to17_3, b17_3to18_3, b18_3to19_3, b19_3to20_3, b20_3to21_3, b21_3to22_3, b22_3to23_3, b23_3to24_3, b24_3to25_3, b25_3to26_3, b26_3to27_3, b27_3to28_3, b28_3to29_3, b29_3to30_3, b30_3to31_3, b31_3to32_3;
wire [`DWIDTH-1:0] b0_4to1_4, b1_4to2_4, b2_4to3_4, b3_4to4_4, b4_4to5_4, b5_4to6_4, b6_4to7_4, b7_4to8_4, b8_4to9_4, b9_4to10_4, b10_4to11_4, b11_4to12_4, b12_4to13_4, b13_4to14_4, b14_4to15_4, b15_4to16_4, b16_4to17_4, b17_4to18_4, b18_4to19_4, b19_4to20_4, b20_4to21_4, b21_4to22_4, b22_4to23_4, b23_4to24_4, b24_4to25_4, b25_4to26_4, b26_4to27_4, b27_4to28_4, b28_4to29_4, b29_4to30_4, b30_4to31_4, b31_4to32_4;
wire [`DWIDTH-1:0] b0_5to1_5, b1_5to2_5, b2_5to3_5, b3_5to4_5, b4_5to5_5, b5_5to6_5, b6_5to7_5, b7_5to8_5, b8_5to9_5, b9_5to10_5, b10_5to11_5, b11_5to12_5, b12_5to13_5, b13_5to14_5, b14_5to15_5, b15_5to16_5, b16_5to17_5, b17_5to18_5, b18_5to19_5, b19_5to20_5, b20_5to21_5, b21_5to22_5, b22_5to23_5, b23_5to24_5, b24_5to25_5, b25_5to26_5, b26_5to27_5, b27_5to28_5, b28_5to29_5, b29_5to30_5, b30_5to31_5, b31_5to32_5;
wire [`DWIDTH-1:0] b0_6to1_6, b1_6to2_6, b2_6to3_6, b3_6to4_6, b4_6to5_6, b5_6to6_6, b6_6to7_6, b7_6to8_6, b8_6to9_6, b9_6to10_6, b10_6to11_6, b11_6to12_6, b12_6to13_6, b13_6to14_6, b14_6to15_6, b15_6to16_6, b16_6to17_6, b17_6to18_6, b18_6to19_6, b19_6to20_6, b20_6to21_6, b21_6to22_6, b22_6to23_6, b23_6to24_6, b24_6to25_6, b25_6to26_6, b26_6to27_6, b27_6to28_6, b28_6to29_6, b29_6to30_6, b30_6to31_6, b31_6to32_6;
wire [`DWIDTH-1:0] b0_7to1_7, b1_7to2_7, b2_7to3_7, b3_7to4_7, b4_7to5_7, b5_7to6_7, b6_7to7_7, b7_7to8_7, b8_7to9_7, b9_7to10_7, b10_7to11_7, b11_7to12_7, b12_7to13_7, b13_7to14_7, b14_7to15_7, b15_7to16_7, b16_7to17_7, b17_7to18_7, b18_7to19_7, b19_7to20_7, b20_7to21_7, b21_7to22_7, b22_7to23_7, b23_7to24_7, b24_7to25_7, b25_7to26_7, b26_7to27_7, b27_7to28_7, b28_7to29_7, b29_7to30_7, b30_7to31_7, b31_7to32_7;
wire [`DWIDTH-1:0] b0_8to1_8, b1_8to2_8, b2_8to3_8, b3_8to4_8, b4_8to5_8, b5_8to6_8, b6_8to7_8, b7_8to8_8, b8_8to9_8, b9_8to10_8, b10_8to11_8, b11_8to12_8, b12_8to13_8, b13_8to14_8, b14_8to15_8, b15_8to16_8, b16_8to17_8, b17_8to18_8, b18_8to19_8, b19_8to20_8, b20_8to21_8, b21_8to22_8, b22_8to23_8, b23_8to24_8, b24_8to25_8, b25_8to26_8, b26_8to27_8, b27_8to28_8, b28_8to29_8, b29_8to30_8, b30_8to31_8, b31_8to32_8;
wire [`DWIDTH-1:0] b0_9to1_9, b1_9to2_9, b2_9to3_9, b3_9to4_9, b4_9to5_9, b5_9to6_9, b6_9to7_9, b7_9to8_9, b8_9to9_9, b9_9to10_9, b10_9to11_9, b11_9to12_9, b12_9to13_9, b13_9to14_9, b14_9to15_9, b15_9to16_9, b16_9to17_9, b17_9to18_9, b18_9to19_9, b19_9to20_9, b20_9to21_9, b21_9to22_9, b22_9to23_9, b23_9to24_9, b24_9to25_9, b25_9to26_9, b26_9to27_9, b27_9to28_9, b28_9to29_9, b29_9to30_9, b30_9to31_9, b31_9to32_9;
wire [`DWIDTH-1:0] b0_10to1_10, b1_10to2_10, b2_10to3_10, b3_10to4_10, b4_10to5_10, b5_10to6_10, b6_10to7_10, b7_10to8_10, b8_10to9_10, b9_10to10_10, b10_10to11_10, b11_10to12_10, b12_10to13_10, b13_10to14_10, b14_10to15_10, b15_10to16_10, b16_10to17_10, b17_10to18_10, b18_10to19_10, b19_10to20_10, b20_10to21_10, b21_10to22_10, b22_10to23_10, b23_10to24_10, b24_10to25_10, b25_10to26_10, b26_10to27_10, b27_10to28_10, b28_10to29_10, b29_10to30_10, b30_10to31_10, b31_10to32_10;
wire [`DWIDTH-1:0] b0_11to1_11, b1_11to2_11, b2_11to3_11, b3_11to4_11, b4_11to5_11, b5_11to6_11, b6_11to7_11, b7_11to8_11, b8_11to9_11, b9_11to10_11, b10_11to11_11, b11_11to12_11, b12_11to13_11, b13_11to14_11, b14_11to15_11, b15_11to16_11, b16_11to17_11, b17_11to18_11, b18_11to19_11, b19_11to20_11, b20_11to21_11, b21_11to22_11, b22_11to23_11, b23_11to24_11, b24_11to25_11, b25_11to26_11, b26_11to27_11, b27_11to28_11, b28_11to29_11, b29_11to30_11, b30_11to31_11, b31_11to32_11;
wire [`DWIDTH-1:0] b0_12to1_12, b1_12to2_12, b2_12to3_12, b3_12to4_12, b4_12to5_12, b5_12to6_12, b6_12to7_12, b7_12to8_12, b8_12to9_12, b9_12to10_12, b10_12to11_12, b11_12to12_12, b12_12to13_12, b13_12to14_12, b14_12to15_12, b15_12to16_12, b16_12to17_12, b17_12to18_12, b18_12to19_12, b19_12to20_12, b20_12to21_12, b21_12to22_12, b22_12to23_12, b23_12to24_12, b24_12to25_12, b25_12to26_12, b26_12to27_12, b27_12to28_12, b28_12to29_12, b29_12to30_12, b30_12to31_12, b31_12to32_12;
wire [`DWIDTH-1:0] b0_13to1_13, b1_13to2_13, b2_13to3_13, b3_13to4_13, b4_13to5_13, b5_13to6_13, b6_13to7_13, b7_13to8_13, b8_13to9_13, b9_13to10_13, b10_13to11_13, b11_13to12_13, b12_13to13_13, b13_13to14_13, b14_13to15_13, b15_13to16_13, b16_13to17_13, b17_13to18_13, b18_13to19_13, b19_13to20_13, b20_13to21_13, b21_13to22_13, b22_13to23_13, b23_13to24_13, b24_13to25_13, b25_13to26_13, b26_13to27_13, b27_13to28_13, b28_13to29_13, b29_13to30_13, b30_13to31_13, b31_13to32_13;
wire [`DWIDTH-1:0] b0_14to1_14, b1_14to2_14, b2_14to3_14, b3_14to4_14, b4_14to5_14, b5_14to6_14, b6_14to7_14, b7_14to8_14, b8_14to9_14, b9_14to10_14, b10_14to11_14, b11_14to12_14, b12_14to13_14, b13_14to14_14, b14_14to15_14, b15_14to16_14, b16_14to17_14, b17_14to18_14, b18_14to19_14, b19_14to20_14, b20_14to21_14, b21_14to22_14, b22_14to23_14, b23_14to24_14, b24_14to25_14, b25_14to26_14, b26_14to27_14, b27_14to28_14, b28_14to29_14, b29_14to30_14, b30_14to31_14, b31_14to32_14;
wire [`DWIDTH-1:0] b0_15to1_15, b1_15to2_15, b2_15to3_15, b3_15to4_15, b4_15to5_15, b5_15to6_15, b6_15to7_15, b7_15to8_15, b8_15to9_15, b9_15to10_15, b10_15to11_15, b11_15to12_15, b12_15to13_15, b13_15to14_15, b14_15to15_15, b15_15to16_15, b16_15to17_15, b17_15to18_15, b18_15to19_15, b19_15to20_15, b20_15to21_15, b21_15to22_15, b22_15to23_15, b23_15to24_15, b24_15to25_15, b25_15to26_15, b26_15to27_15, b27_15to28_15, b28_15to29_15, b29_15to30_15, b30_15to31_15, b31_15to32_15;
wire [`DWIDTH-1:0] b0_16to1_16, b1_16to2_16, b2_16to3_16, b3_16to4_16, b4_16to5_16, b5_16to6_16, b6_16to7_16, b7_16to8_16, b8_16to9_16, b9_16to10_16, b10_16to11_16, b11_16to12_16, b12_16to13_16, b13_16to14_16, b14_16to15_16, b15_16to16_16, b16_16to17_16, b17_16to18_16, b18_16to19_16, b19_16to20_16, b20_16to21_16, b21_16to22_16, b22_16to23_16, b23_16to24_16, b24_16to25_16, b25_16to26_16, b26_16to27_16, b27_16to28_16, b28_16to29_16, b29_16to30_16, b30_16to31_16, b31_16to32_16;
wire [`DWIDTH-1:0] b0_17to1_17, b1_17to2_17, b2_17to3_17, b3_17to4_17, b4_17to5_17, b5_17to6_17, b6_17to7_17, b7_17to8_17, b8_17to9_17, b9_17to10_17, b10_17to11_17, b11_17to12_17, b12_17to13_17, b13_17to14_17, b14_17to15_17, b15_17to16_17, b16_17to17_17, b17_17to18_17, b18_17to19_17, b19_17to20_17, b20_17to21_17, b21_17to22_17, b22_17to23_17, b23_17to24_17, b24_17to25_17, b25_17to26_17, b26_17to27_17, b27_17to28_17, b28_17to29_17, b29_17to30_17, b30_17to31_17, b31_17to32_17;
wire [`DWIDTH-1:0] b0_18to1_18, b1_18to2_18, b2_18to3_18, b3_18to4_18, b4_18to5_18, b5_18to6_18, b6_18to7_18, b7_18to8_18, b8_18to9_18, b9_18to10_18, b10_18to11_18, b11_18to12_18, b12_18to13_18, b13_18to14_18, b14_18to15_18, b15_18to16_18, b16_18to17_18, b17_18to18_18, b18_18to19_18, b19_18to20_18, b20_18to21_18, b21_18to22_18, b22_18to23_18, b23_18to24_18, b24_18to25_18, b25_18to26_18, b26_18to27_18, b27_18to28_18, b28_18to29_18, b29_18to30_18, b30_18to31_18, b31_18to32_18;
wire [`DWIDTH-1:0] b0_19to1_19, b1_19to2_19, b2_19to3_19, b3_19to4_19, b4_19to5_19, b5_19to6_19, b6_19to7_19, b7_19to8_19, b8_19to9_19, b9_19to10_19, b10_19to11_19, b11_19to12_19, b12_19to13_19, b13_19to14_19, b14_19to15_19, b15_19to16_19, b16_19to17_19, b17_19to18_19, b18_19to19_19, b19_19to20_19, b20_19to21_19, b21_19to22_19, b22_19to23_19, b23_19to24_19, b24_19to25_19, b25_19to26_19, b26_19to27_19, b27_19to28_19, b28_19to29_19, b29_19to30_19, b30_19to31_19, b31_19to32_19;
wire [`DWIDTH-1:0] b0_20to1_20, b1_20to2_20, b2_20to3_20, b3_20to4_20, b4_20to5_20, b5_20to6_20, b6_20to7_20, b7_20to8_20, b8_20to9_20, b9_20to10_20, b10_20to11_20, b11_20to12_20, b12_20to13_20, b13_20to14_20, b14_20to15_20, b15_20to16_20, b16_20to17_20, b17_20to18_20, b18_20to19_20, b19_20to20_20, b20_20to21_20, b21_20to22_20, b22_20to23_20, b23_20to24_20, b24_20to25_20, b25_20to26_20, b26_20to27_20, b27_20to28_20, b28_20to29_20, b29_20to30_20, b30_20to31_20, b31_20to32_20;
wire [`DWIDTH-1:0] b0_21to1_21, b1_21to2_21, b2_21to3_21, b3_21to4_21, b4_21to5_21, b5_21to6_21, b6_21to7_21, b7_21to8_21, b8_21to9_21, b9_21to10_21, b10_21to11_21, b11_21to12_21, b12_21to13_21, b13_21to14_21, b14_21to15_21, b15_21to16_21, b16_21to17_21, b17_21to18_21, b18_21to19_21, b19_21to20_21, b20_21to21_21, b21_21to22_21, b22_21to23_21, b23_21to24_21, b24_21to25_21, b25_21to26_21, b26_21to27_21, b27_21to28_21, b28_21to29_21, b29_21to30_21, b30_21to31_21, b31_21to32_21;
wire [`DWIDTH-1:0] b0_22to1_22, b1_22to2_22, b2_22to3_22, b3_22to4_22, b4_22to5_22, b5_22to6_22, b6_22to7_22, b7_22to8_22, b8_22to9_22, b9_22to10_22, b10_22to11_22, b11_22to12_22, b12_22to13_22, b13_22to14_22, b14_22to15_22, b15_22to16_22, b16_22to17_22, b17_22to18_22, b18_22to19_22, b19_22to20_22, b20_22to21_22, b21_22to22_22, b22_22to23_22, b23_22to24_22, b24_22to25_22, b25_22to26_22, b26_22to27_22, b27_22to28_22, b28_22to29_22, b29_22to30_22, b30_22to31_22, b31_22to32_22;
wire [`DWIDTH-1:0] b0_23to1_23, b1_23to2_23, b2_23to3_23, b3_23to4_23, b4_23to5_23, b5_23to6_23, b6_23to7_23, b7_23to8_23, b8_23to9_23, b9_23to10_23, b10_23to11_23, b11_23to12_23, b12_23to13_23, b13_23to14_23, b14_23to15_23, b15_23to16_23, b16_23to17_23, b17_23to18_23, b18_23to19_23, b19_23to20_23, b20_23to21_23, b21_23to22_23, b22_23to23_23, b23_23to24_23, b24_23to25_23, b25_23to26_23, b26_23to27_23, b27_23to28_23, b28_23to29_23, b29_23to30_23, b30_23to31_23, b31_23to32_23;
wire [`DWIDTH-1:0] b0_24to1_24, b1_24to2_24, b2_24to3_24, b3_24to4_24, b4_24to5_24, b5_24to6_24, b6_24to7_24, b7_24to8_24, b8_24to9_24, b9_24to10_24, b10_24to11_24, b11_24to12_24, b12_24to13_24, b13_24to14_24, b14_24to15_24, b15_24to16_24, b16_24to17_24, b17_24to18_24, b18_24to19_24, b19_24to20_24, b20_24to21_24, b21_24to22_24, b22_24to23_24, b23_24to24_24, b24_24to25_24, b25_24to26_24, b26_24to27_24, b27_24to28_24, b28_24to29_24, b29_24to30_24, b30_24to31_24, b31_24to32_24;
wire [`DWIDTH-1:0] b0_25to1_25, b1_25to2_25, b2_25to3_25, b3_25to4_25, b4_25to5_25, b5_25to6_25, b6_25to7_25, b7_25to8_25, b8_25to9_25, b9_25to10_25, b10_25to11_25, b11_25to12_25, b12_25to13_25, b13_25to14_25, b14_25to15_25, b15_25to16_25, b16_25to17_25, b17_25to18_25, b18_25to19_25, b19_25to20_25, b20_25to21_25, b21_25to22_25, b22_25to23_25, b23_25to24_25, b24_25to25_25, b25_25to26_25, b26_25to27_25, b27_25to28_25, b28_25to29_25, b29_25to30_25, b30_25to31_25, b31_25to32_25;
wire [`DWIDTH-1:0] b0_26to1_26, b1_26to2_26, b2_26to3_26, b3_26to4_26, b4_26to5_26, b5_26to6_26, b6_26to7_26, b7_26to8_26, b8_26to9_26, b9_26to10_26, b10_26to11_26, b11_26to12_26, b12_26to13_26, b13_26to14_26, b14_26to15_26, b15_26to16_26, b16_26to17_26, b17_26to18_26, b18_26to19_26, b19_26to20_26, b20_26to21_26, b21_26to22_26, b22_26to23_26, b23_26to24_26, b24_26to25_26, b25_26to26_26, b26_26to27_26, b27_26to28_26, b28_26to29_26, b29_26to30_26, b30_26to31_26, b31_26to32_26;
wire [`DWIDTH-1:0] b0_27to1_27, b1_27to2_27, b2_27to3_27, b3_27to4_27, b4_27to5_27, b5_27to6_27, b6_27to7_27, b7_27to8_27, b8_27to9_27, b9_27to10_27, b10_27to11_27, b11_27to12_27, b12_27to13_27, b13_27to14_27, b14_27to15_27, b15_27to16_27, b16_27to17_27, b17_27to18_27, b18_27to19_27, b19_27to20_27, b20_27to21_27, b21_27to22_27, b22_27to23_27, b23_27to24_27, b24_27to25_27, b25_27to26_27, b26_27to27_27, b27_27to28_27, b28_27to29_27, b29_27to30_27, b30_27to31_27, b31_27to32_27;
wire [`DWIDTH-1:0] b0_28to1_28, b1_28to2_28, b2_28to3_28, b3_28to4_28, b4_28to5_28, b5_28to6_28, b6_28to7_28, b7_28to8_28, b8_28to9_28, b9_28to10_28, b10_28to11_28, b11_28to12_28, b12_28to13_28, b13_28to14_28, b14_28to15_28, b15_28to16_28, b16_28to17_28, b17_28to18_28, b18_28to19_28, b19_28to20_28, b20_28to21_28, b21_28to22_28, b22_28to23_28, b23_28to24_28, b24_28to25_28, b25_28to26_28, b26_28to27_28, b27_28to28_28, b28_28to29_28, b29_28to30_28, b30_28to31_28, b31_28to32_28;
wire [`DWIDTH-1:0] b0_29to1_29, b1_29to2_29, b2_29to3_29, b3_29to4_29, b4_29to5_29, b5_29to6_29, b6_29to7_29, b7_29to8_29, b8_29to9_29, b9_29to10_29, b10_29to11_29, b11_29to12_29, b12_29to13_29, b13_29to14_29, b14_29to15_29, b15_29to16_29, b16_29to17_29, b17_29to18_29, b18_29to19_29, b19_29to20_29, b20_29to21_29, b21_29to22_29, b22_29to23_29, b23_29to24_29, b24_29to25_29, b25_29to26_29, b26_29to27_29, b27_29to28_29, b28_29to29_29, b29_29to30_29, b30_29to31_29, b31_29to32_29;
wire [`DWIDTH-1:0] b0_30to1_30, b1_30to2_30, b2_30to3_30, b3_30to4_30, b4_30to5_30, b5_30to6_30, b6_30to7_30, b7_30to8_30, b8_30to9_30, b9_30to10_30, b10_30to11_30, b11_30to12_30, b12_30to13_30, b13_30to14_30, b14_30to15_30, b15_30to16_30, b16_30to17_30, b17_30to18_30, b18_30to19_30, b19_30to20_30, b20_30to21_30, b21_30to22_30, b22_30to23_30, b23_30to24_30, b24_30to25_30, b25_30to26_30, b26_30to27_30, b27_30to28_30, b28_30to29_30, b29_30to30_30, b30_30to31_30, b31_30to32_30;
wire [`DWIDTH-1:0] b0_31to1_31, b1_31to2_31, b2_31to3_31, b3_31to4_31, b4_31to5_31, b5_31to6_31, b6_31to7_31, b7_31to8_31, b8_31to9_31, b9_31to10_31, b10_31to11_31, b11_31to12_31, b12_31to13_31, b13_31to14_31, b14_31to15_31, b15_31to16_31, b16_31to17_31, b17_31to18_31, b18_31to19_31, b19_31to20_31, b20_31to21_31, b21_31to22_31, b22_31to23_31, b23_31to24_31, b24_31to25_31, b25_31to26_31, b26_31to27_31, b27_31to28_31, b28_31to29_31, b29_31to30_31, b30_31to31_31, b31_31to32_31;

//////////////////////////////////////////////////////////////////////////
// Instantiations of the actual PEs
//////////////////////////////////////////////////////////////////////////
//For larger matmul, more PEs will be needed
wire effective_rst;
assign effective_rst = reset | pe_reset;

processing_element pe0_0(.reset(effective_rst), .clk(clk),  .in_a(a0),      .in_b(b0),  .out_a(a0_0to0_1), .out_b(b0_0to1_0), .out_c(matrixC0_0));
processing_element pe0_1(.reset(effective_rst), .clk(clk),  .in_a(a0_0to0_1), .in_b(b1),  .out_a(a0_1to0_2), .out_b(b0_1to1_1), .out_c(matrixC0_1));
processing_element pe0_2(.reset(effective_rst), .clk(clk),  .in_a(a0_1to0_2), .in_b(b2),  .out_a(a0_2to0_3), .out_b(b0_2to1_2), .out_c(matrixC0_2));
processing_element pe0_3(.reset(effective_rst), .clk(clk),  .in_a(a0_2to0_3), .in_b(b3),  .out_a(a0_3to0_4), .out_b(b0_3to1_3), .out_c(matrixC0_3));
processing_element pe0_4(.reset(effective_rst), .clk(clk),  .in_a(a0_3to0_4), .in_b(b4),  .out_a(a0_4to0_5), .out_b(b0_4to1_4), .out_c(matrixC0_4));
processing_element pe0_5(.reset(effective_rst), .clk(clk),  .in_a(a0_4to0_5), .in_b(b5),  .out_a(a0_5to0_6), .out_b(b0_5to1_5), .out_c(matrixC0_5));
processing_element pe0_6(.reset(effective_rst), .clk(clk),  .in_a(a0_5to0_6), .in_b(b6),  .out_a(a0_6to0_7), .out_b(b0_6to1_6), .out_c(matrixC0_6));
processing_element pe0_7(.reset(effective_rst), .clk(clk),  .in_a(a0_6to0_7), .in_b(b7),  .out_a(a0_7to0_8), .out_b(b0_7to1_7), .out_c(matrixC0_7));
processing_element pe0_8(.reset(effective_rst), .clk(clk),  .in_a(a0_7to0_8), .in_b(b8),  .out_a(a0_8to0_9), .out_b(b0_8to1_8), .out_c(matrixC0_8));
processing_element pe0_9(.reset(effective_rst), .clk(clk),  .in_a(a0_8to0_9), .in_b(b9),  .out_a(a0_9to0_10), .out_b(b0_9to1_9), .out_c(matrixC0_9));
processing_element pe0_10(.reset(effective_rst), .clk(clk),  .in_a(a0_9to0_10), .in_b(b10),  .out_a(a0_10to0_11), .out_b(b0_10to1_10), .out_c(matrixC0_10));
processing_element pe0_11(.reset(effective_rst), .clk(clk),  .in_a(a0_10to0_11), .in_b(b11),  .out_a(a0_11to0_12), .out_b(b0_11to1_11), .out_c(matrixC0_11));
processing_element pe0_12(.reset(effective_rst), .clk(clk),  .in_a(a0_11to0_12), .in_b(b12),  .out_a(a0_12to0_13), .out_b(b0_12to1_12), .out_c(matrixC0_12));
processing_element pe0_13(.reset(effective_rst), .clk(clk),  .in_a(a0_12to0_13), .in_b(b13),  .out_a(a0_13to0_14), .out_b(b0_13to1_13), .out_c(matrixC0_13));
processing_element pe0_14(.reset(effective_rst), .clk(clk),  .in_a(a0_13to0_14), .in_b(b14),  .out_a(a0_14to0_15), .out_b(b0_14to1_14), .out_c(matrixC0_14));
processing_element pe0_15(.reset(effective_rst), .clk(clk),  .in_a(a0_14to0_15), .in_b(b15),  .out_a(a0_15to0_16), .out_b(b0_15to1_15), .out_c(matrixC0_15));
processing_element pe0_16(.reset(effective_rst), .clk(clk),  .in_a(a0_15to0_16), .in_b(b16),  .out_a(a0_16to0_17), .out_b(b0_16to1_16), .out_c(matrixC0_16));
processing_element pe0_17(.reset(effective_rst), .clk(clk),  .in_a(a0_16to0_17), .in_b(b17),  .out_a(a0_17to0_18), .out_b(b0_17to1_17), .out_c(matrixC0_17));
processing_element pe0_18(.reset(effective_rst), .clk(clk),  .in_a(a0_17to0_18), .in_b(b18),  .out_a(a0_18to0_19), .out_b(b0_18to1_18), .out_c(matrixC0_18));
processing_element pe0_19(.reset(effective_rst), .clk(clk),  .in_a(a0_18to0_19), .in_b(b19),  .out_a(a0_19to0_20), .out_b(b0_19to1_19), .out_c(matrixC0_19));
processing_element pe0_20(.reset(effective_rst), .clk(clk),  .in_a(a0_19to0_20), .in_b(b20),  .out_a(a0_20to0_21), .out_b(b0_20to1_20), .out_c(matrixC0_20));
processing_element pe0_21(.reset(effective_rst), .clk(clk),  .in_a(a0_20to0_21), .in_b(b21),  .out_a(a0_21to0_22), .out_b(b0_21to1_21), .out_c(matrixC0_21));
processing_element pe0_22(.reset(effective_rst), .clk(clk),  .in_a(a0_21to0_22), .in_b(b22),  .out_a(a0_22to0_23), .out_b(b0_22to1_22), .out_c(matrixC0_22));
processing_element pe0_23(.reset(effective_rst), .clk(clk),  .in_a(a0_22to0_23), .in_b(b23),  .out_a(a0_23to0_24), .out_b(b0_23to1_23), .out_c(matrixC0_23));
processing_element pe0_24(.reset(effective_rst), .clk(clk),  .in_a(a0_23to0_24), .in_b(b24),  .out_a(a0_24to0_25), .out_b(b0_24to1_24), .out_c(matrixC0_24));
processing_element pe0_25(.reset(effective_rst), .clk(clk),  .in_a(a0_24to0_25), .in_b(b25),  .out_a(a0_25to0_26), .out_b(b0_25to1_25), .out_c(matrixC0_25));
processing_element pe0_26(.reset(effective_rst), .clk(clk),  .in_a(a0_25to0_26), .in_b(b26),  .out_a(a0_26to0_27), .out_b(b0_26to1_26), .out_c(matrixC0_26));
processing_element pe0_27(.reset(effective_rst), .clk(clk),  .in_a(a0_26to0_27), .in_b(b27),  .out_a(a0_27to0_28), .out_b(b0_27to1_27), .out_c(matrixC0_27));
processing_element pe0_28(.reset(effective_rst), .clk(clk),  .in_a(a0_27to0_28), .in_b(b28),  .out_a(a0_28to0_29), .out_b(b0_28to1_28), .out_c(matrixC0_28));
processing_element pe0_29(.reset(effective_rst), .clk(clk),  .in_a(a0_28to0_29), .in_b(b29),  .out_a(a0_29to0_30), .out_b(b0_29to1_29), .out_c(matrixC0_29));
processing_element pe0_30(.reset(effective_rst), .clk(clk),  .in_a(a0_29to0_30), .in_b(b30),  .out_a(a0_30to0_31), .out_b(b0_30to1_30), .out_c(matrixC0_30));
processing_element pe0_31(.reset(effective_rst), .clk(clk),  .in_a(a0_30to0_31), .in_b(b31),  .out_a(a0_31to0_32), .out_b(b0_31to1_31), .out_c(matrixC0_31));

processing_element pe1_0(.reset(effective_rst), .clk(clk),  .in_a(a1), .in_b(b0_0to1_0),  .out_a(a1_0to1_1), .out_b(b1_0to2_0), .out_c(matrixC1_0));
processing_element pe2_0(.reset(effective_rst), .clk(clk),  .in_a(a2), .in_b(b1_0to2_0),  .out_a(a2_0to2_1), .out_b(b2_0to3_0), .out_c(matrixC2_0));
processing_element pe3_0(.reset(effective_rst), .clk(clk),  .in_a(a3), .in_b(b2_0to3_0),  .out_a(a3_0to3_1), .out_b(b3_0to4_0), .out_c(matrixC3_0));
processing_element pe4_0(.reset(effective_rst), .clk(clk),  .in_a(a4), .in_b(b3_0to4_0),  .out_a(a4_0to4_1), .out_b(b4_0to5_0), .out_c(matrixC4_0));
processing_element pe5_0(.reset(effective_rst), .clk(clk),  .in_a(a5), .in_b(b4_0to5_0),  .out_a(a5_0to5_1), .out_b(b5_0to6_0), .out_c(matrixC5_0));
processing_element pe6_0(.reset(effective_rst), .clk(clk),  .in_a(a6), .in_b(b5_0to6_0),  .out_a(a6_0to6_1), .out_b(b6_0to7_0), .out_c(matrixC6_0));
processing_element pe7_0(.reset(effective_rst), .clk(clk),  .in_a(a7), .in_b(b6_0to7_0),  .out_a(a7_0to7_1), .out_b(b7_0to8_0), .out_c(matrixC7_0));
processing_element pe8_0(.reset(effective_rst), .clk(clk),  .in_a(a8), .in_b(b7_0to8_0),  .out_a(a8_0to8_1), .out_b(b8_0to9_0), .out_c(matrixC8_0));
processing_element pe9_0(.reset(effective_rst), .clk(clk),  .in_a(a9), .in_b(b8_0to9_0),  .out_a(a9_0to9_1), .out_b(b9_0to10_0), .out_c(matrixC9_0));
processing_element pe10_0(.reset(effective_rst), .clk(clk),  .in_a(a10), .in_b(b9_0to10_0),  .out_a(a10_0to10_1), .out_b(b10_0to11_0), .out_c(matrixC10_0));
processing_element pe11_0(.reset(effective_rst), .clk(clk),  .in_a(a11), .in_b(b10_0to11_0),  .out_a(a11_0to11_1), .out_b(b11_0to12_0), .out_c(matrixC11_0));
processing_element pe12_0(.reset(effective_rst), .clk(clk),  .in_a(a12), .in_b(b11_0to12_0),  .out_a(a12_0to12_1), .out_b(b12_0to13_0), .out_c(matrixC12_0));
processing_element pe13_0(.reset(effective_rst), .clk(clk),  .in_a(a13), .in_b(b12_0to13_0),  .out_a(a13_0to13_1), .out_b(b13_0to14_0), .out_c(matrixC13_0));
processing_element pe14_0(.reset(effective_rst), .clk(clk),  .in_a(a14), .in_b(b13_0to14_0),  .out_a(a14_0to14_1), .out_b(b14_0to15_0), .out_c(matrixC14_0));
processing_element pe15_0(.reset(effective_rst), .clk(clk),  .in_a(a15), .in_b(b14_0to15_0),  .out_a(a15_0to15_1), .out_b(b15_0to16_0), .out_c(matrixC15_0));
processing_element pe16_0(.reset(effective_rst), .clk(clk),  .in_a(a16), .in_b(b15_0to16_0),  .out_a(a16_0to16_1), .out_b(b16_0to17_0), .out_c(matrixC16_0));
processing_element pe17_0(.reset(effective_rst), .clk(clk),  .in_a(a17), .in_b(b16_0to17_0),  .out_a(a17_0to17_1), .out_b(b17_0to18_0), .out_c(matrixC17_0));
processing_element pe18_0(.reset(effective_rst), .clk(clk),  .in_a(a18), .in_b(b17_0to18_0),  .out_a(a18_0to18_1), .out_b(b18_0to19_0), .out_c(matrixC18_0));
processing_element pe19_0(.reset(effective_rst), .clk(clk),  .in_a(a19), .in_b(b18_0to19_0),  .out_a(a19_0to19_1), .out_b(b19_0to20_0), .out_c(matrixC19_0));
processing_element pe20_0(.reset(effective_rst), .clk(clk),  .in_a(a20), .in_b(b19_0to20_0),  .out_a(a20_0to20_1), .out_b(b20_0to21_0), .out_c(matrixC20_0));
processing_element pe21_0(.reset(effective_rst), .clk(clk),  .in_a(a21), .in_b(b20_0to21_0),  .out_a(a21_0to21_1), .out_b(b21_0to22_0), .out_c(matrixC21_0));
processing_element pe22_0(.reset(effective_rst), .clk(clk),  .in_a(a22), .in_b(b21_0to22_0),  .out_a(a22_0to22_1), .out_b(b22_0to23_0), .out_c(matrixC22_0));
processing_element pe23_0(.reset(effective_rst), .clk(clk),  .in_a(a23), .in_b(b22_0to23_0),  .out_a(a23_0to23_1), .out_b(b23_0to24_0), .out_c(matrixC23_0));
processing_element pe24_0(.reset(effective_rst), .clk(clk),  .in_a(a24), .in_b(b23_0to24_0),  .out_a(a24_0to24_1), .out_b(b24_0to25_0), .out_c(matrixC24_0));
processing_element pe25_0(.reset(effective_rst), .clk(clk),  .in_a(a25), .in_b(b24_0to25_0),  .out_a(a25_0to25_1), .out_b(b25_0to26_0), .out_c(matrixC25_0));
processing_element pe26_0(.reset(effective_rst), .clk(clk),  .in_a(a26), .in_b(b25_0to26_0),  .out_a(a26_0to26_1), .out_b(b26_0to27_0), .out_c(matrixC26_0));
processing_element pe27_0(.reset(effective_rst), .clk(clk),  .in_a(a27), .in_b(b26_0to27_0),  .out_a(a27_0to27_1), .out_b(b27_0to28_0), .out_c(matrixC27_0));
processing_element pe28_0(.reset(effective_rst), .clk(clk),  .in_a(a28), .in_b(b27_0to28_0),  .out_a(a28_0to28_1), .out_b(b28_0to29_0), .out_c(matrixC28_0));
processing_element pe29_0(.reset(effective_rst), .clk(clk),  .in_a(a29), .in_b(b28_0to29_0),  .out_a(a29_0to29_1), .out_b(b29_0to30_0), .out_c(matrixC29_0));
processing_element pe30_0(.reset(effective_rst), .clk(clk),  .in_a(a30), .in_b(b29_0to30_0),  .out_a(a30_0to30_1), .out_b(b30_0to31_0), .out_c(matrixC30_0));
processing_element pe31_0(.reset(effective_rst), .clk(clk),  .in_a(a31), .in_b(b30_0to31_0),  .out_a(a31_0to31_1), .out_b(b31_0to32_0), .out_c(matrixC31_0));

processing_element pe1_1(.reset(effective_rst), .clk(clk),  .in_a(a1_0to1_1), .in_b(b0_1to1_1),  .out_a(a1_1to1_2), .out_b(b1_1to2_1), .out_c(matrixC1_1));
processing_element pe1_2(.reset(effective_rst), .clk(clk),  .in_a(a1_1to1_2), .in_b(b0_2to1_2),  .out_a(a1_2to1_3), .out_b(b1_2to2_2), .out_c(matrixC1_2));
processing_element pe1_3(.reset(effective_rst), .clk(clk),  .in_a(a1_2to1_3), .in_b(b0_3to1_3),  .out_a(a1_3to1_4), .out_b(b1_3to2_3), .out_c(matrixC1_3));
processing_element pe1_4(.reset(effective_rst), .clk(clk),  .in_a(a1_3to1_4), .in_b(b0_4to1_4),  .out_a(a1_4to1_5), .out_b(b1_4to2_4), .out_c(matrixC1_4));
processing_element pe1_5(.reset(effective_rst), .clk(clk),  .in_a(a1_4to1_5), .in_b(b0_5to1_5),  .out_a(a1_5to1_6), .out_b(b1_5to2_5), .out_c(matrixC1_5));
processing_element pe1_6(.reset(effective_rst), .clk(clk),  .in_a(a1_5to1_6), .in_b(b0_6to1_6),  .out_a(a1_6to1_7), .out_b(b1_6to2_6), .out_c(matrixC1_6));
processing_element pe1_7(.reset(effective_rst), .clk(clk),  .in_a(a1_6to1_7), .in_b(b0_7to1_7),  .out_a(a1_7to1_8), .out_b(b1_7to2_7), .out_c(matrixC1_7));
processing_element pe1_8(.reset(effective_rst), .clk(clk),  .in_a(a1_7to1_8), .in_b(b0_8to1_8),  .out_a(a1_8to1_9), .out_b(b1_8to2_8), .out_c(matrixC1_8));
processing_element pe1_9(.reset(effective_rst), .clk(clk),  .in_a(a1_8to1_9), .in_b(b0_9to1_9),  .out_a(a1_9to1_10), .out_b(b1_9to2_9), .out_c(matrixC1_9));
processing_element pe1_10(.reset(effective_rst), .clk(clk),  .in_a(a1_9to1_10), .in_b(b0_10to1_10),  .out_a(a1_10to1_11), .out_b(b1_10to2_10), .out_c(matrixC1_10));
processing_element pe1_11(.reset(effective_rst), .clk(clk),  .in_a(a1_10to1_11), .in_b(b0_11to1_11),  .out_a(a1_11to1_12), .out_b(b1_11to2_11), .out_c(matrixC1_11));
processing_element pe1_12(.reset(effective_rst), .clk(clk),  .in_a(a1_11to1_12), .in_b(b0_12to1_12),  .out_a(a1_12to1_13), .out_b(b1_12to2_12), .out_c(matrixC1_12));
processing_element pe1_13(.reset(effective_rst), .clk(clk),  .in_a(a1_12to1_13), .in_b(b0_13to1_13),  .out_a(a1_13to1_14), .out_b(b1_13to2_13), .out_c(matrixC1_13));
processing_element pe1_14(.reset(effective_rst), .clk(clk),  .in_a(a1_13to1_14), .in_b(b0_14to1_14),  .out_a(a1_14to1_15), .out_b(b1_14to2_14), .out_c(matrixC1_14));
processing_element pe1_15(.reset(effective_rst), .clk(clk),  .in_a(a1_14to1_15), .in_b(b0_15to1_15),  .out_a(a1_15to1_16), .out_b(b1_15to2_15), .out_c(matrixC1_15));
processing_element pe1_16(.reset(effective_rst), .clk(clk),  .in_a(a1_15to1_16), .in_b(b0_16to1_16),  .out_a(a1_16to1_17), .out_b(b1_16to2_16), .out_c(matrixC1_16));
processing_element pe1_17(.reset(effective_rst), .clk(clk),  .in_a(a1_16to1_17), .in_b(b0_17to1_17),  .out_a(a1_17to1_18), .out_b(b1_17to2_17), .out_c(matrixC1_17));
processing_element pe1_18(.reset(effective_rst), .clk(clk),  .in_a(a1_17to1_18), .in_b(b0_18to1_18),  .out_a(a1_18to1_19), .out_b(b1_18to2_18), .out_c(matrixC1_18));
processing_element pe1_19(.reset(effective_rst), .clk(clk),  .in_a(a1_18to1_19), .in_b(b0_19to1_19),  .out_a(a1_19to1_20), .out_b(b1_19to2_19), .out_c(matrixC1_19));
processing_element pe1_20(.reset(effective_rst), .clk(clk),  .in_a(a1_19to1_20), .in_b(b0_20to1_20),  .out_a(a1_20to1_21), .out_b(b1_20to2_20), .out_c(matrixC1_20));
processing_element pe1_21(.reset(effective_rst), .clk(clk),  .in_a(a1_20to1_21), .in_b(b0_21to1_21),  .out_a(a1_21to1_22), .out_b(b1_21to2_21), .out_c(matrixC1_21));
processing_element pe1_22(.reset(effective_rst), .clk(clk),  .in_a(a1_21to1_22), .in_b(b0_22to1_22),  .out_a(a1_22to1_23), .out_b(b1_22to2_22), .out_c(matrixC1_22));
processing_element pe1_23(.reset(effective_rst), .clk(clk),  .in_a(a1_22to1_23), .in_b(b0_23to1_23),  .out_a(a1_23to1_24), .out_b(b1_23to2_23), .out_c(matrixC1_23));
processing_element pe1_24(.reset(effective_rst), .clk(clk),  .in_a(a1_23to1_24), .in_b(b0_24to1_24),  .out_a(a1_24to1_25), .out_b(b1_24to2_24), .out_c(matrixC1_24));
processing_element pe1_25(.reset(effective_rst), .clk(clk),  .in_a(a1_24to1_25), .in_b(b0_25to1_25),  .out_a(a1_25to1_26), .out_b(b1_25to2_25), .out_c(matrixC1_25));
processing_element pe1_26(.reset(effective_rst), .clk(clk),  .in_a(a1_25to1_26), .in_b(b0_26to1_26),  .out_a(a1_26to1_27), .out_b(b1_26to2_26), .out_c(matrixC1_26));
processing_element pe1_27(.reset(effective_rst), .clk(clk),  .in_a(a1_26to1_27), .in_b(b0_27to1_27),  .out_a(a1_27to1_28), .out_b(b1_27to2_27), .out_c(matrixC1_27));
processing_element pe1_28(.reset(effective_rst), .clk(clk),  .in_a(a1_27to1_28), .in_b(b0_28to1_28),  .out_a(a1_28to1_29), .out_b(b1_28to2_28), .out_c(matrixC1_28));
processing_element pe1_29(.reset(effective_rst), .clk(clk),  .in_a(a1_28to1_29), .in_b(b0_29to1_29),  .out_a(a1_29to1_30), .out_b(b1_29to2_29), .out_c(matrixC1_29));
processing_element pe1_30(.reset(effective_rst), .clk(clk),  .in_a(a1_29to1_30), .in_b(b0_30to1_30),  .out_a(a1_30to1_31), .out_b(b1_30to2_30), .out_c(matrixC1_30));
processing_element pe1_31(.reset(effective_rst), .clk(clk),  .in_a(a1_30to1_31), .in_b(b0_31to1_31),  .out_a(a1_31to1_32), .out_b(b1_31to2_31), .out_c(matrixC1_31));
processing_element pe2_1(.reset(effective_rst), .clk(clk),  .in_a(a2_0to2_1), .in_b(b1_1to2_1),  .out_a(a2_1to2_2), .out_b(b2_1to3_1), .out_c(matrixC2_1));
processing_element pe2_2(.reset(effective_rst), .clk(clk),  .in_a(a2_1to2_2), .in_b(b1_2to2_2),  .out_a(a2_2to2_3), .out_b(b2_2to3_2), .out_c(matrixC2_2));
processing_element pe2_3(.reset(effective_rst), .clk(clk),  .in_a(a2_2to2_3), .in_b(b1_3to2_3),  .out_a(a2_3to2_4), .out_b(b2_3to3_3), .out_c(matrixC2_3));
processing_element pe2_4(.reset(effective_rst), .clk(clk),  .in_a(a2_3to2_4), .in_b(b1_4to2_4),  .out_a(a2_4to2_5), .out_b(b2_4to3_4), .out_c(matrixC2_4));
processing_element pe2_5(.reset(effective_rst), .clk(clk),  .in_a(a2_4to2_5), .in_b(b1_5to2_5),  .out_a(a2_5to2_6), .out_b(b2_5to3_5), .out_c(matrixC2_5));
processing_element pe2_6(.reset(effective_rst), .clk(clk),  .in_a(a2_5to2_6), .in_b(b1_6to2_6),  .out_a(a2_6to2_7), .out_b(b2_6to3_6), .out_c(matrixC2_6));
processing_element pe2_7(.reset(effective_rst), .clk(clk),  .in_a(a2_6to2_7), .in_b(b1_7to2_7),  .out_a(a2_7to2_8), .out_b(b2_7to3_7), .out_c(matrixC2_7));
processing_element pe2_8(.reset(effective_rst), .clk(clk),  .in_a(a2_7to2_8), .in_b(b1_8to2_8),  .out_a(a2_8to2_9), .out_b(b2_8to3_8), .out_c(matrixC2_8));
processing_element pe2_9(.reset(effective_rst), .clk(clk),  .in_a(a2_8to2_9), .in_b(b1_9to2_9),  .out_a(a2_9to2_10), .out_b(b2_9to3_9), .out_c(matrixC2_9));
processing_element pe2_10(.reset(effective_rst), .clk(clk),  .in_a(a2_9to2_10), .in_b(b1_10to2_10),  .out_a(a2_10to2_11), .out_b(b2_10to3_10), .out_c(matrixC2_10));
processing_element pe2_11(.reset(effective_rst), .clk(clk),  .in_a(a2_10to2_11), .in_b(b1_11to2_11),  .out_a(a2_11to2_12), .out_b(b2_11to3_11), .out_c(matrixC2_11));
processing_element pe2_12(.reset(effective_rst), .clk(clk),  .in_a(a2_11to2_12), .in_b(b1_12to2_12),  .out_a(a2_12to2_13), .out_b(b2_12to3_12), .out_c(matrixC2_12));
processing_element pe2_13(.reset(effective_rst), .clk(clk),  .in_a(a2_12to2_13), .in_b(b1_13to2_13),  .out_a(a2_13to2_14), .out_b(b2_13to3_13), .out_c(matrixC2_13));
processing_element pe2_14(.reset(effective_rst), .clk(clk),  .in_a(a2_13to2_14), .in_b(b1_14to2_14),  .out_a(a2_14to2_15), .out_b(b2_14to3_14), .out_c(matrixC2_14));
processing_element pe2_15(.reset(effective_rst), .clk(clk),  .in_a(a2_14to2_15), .in_b(b1_15to2_15),  .out_a(a2_15to2_16), .out_b(b2_15to3_15), .out_c(matrixC2_15));
processing_element pe2_16(.reset(effective_rst), .clk(clk),  .in_a(a2_15to2_16), .in_b(b1_16to2_16),  .out_a(a2_16to2_17), .out_b(b2_16to3_16), .out_c(matrixC2_16));
processing_element pe2_17(.reset(effective_rst), .clk(clk),  .in_a(a2_16to2_17), .in_b(b1_17to2_17),  .out_a(a2_17to2_18), .out_b(b2_17to3_17), .out_c(matrixC2_17));
processing_element pe2_18(.reset(effective_rst), .clk(clk),  .in_a(a2_17to2_18), .in_b(b1_18to2_18),  .out_a(a2_18to2_19), .out_b(b2_18to3_18), .out_c(matrixC2_18));
processing_element pe2_19(.reset(effective_rst), .clk(clk),  .in_a(a2_18to2_19), .in_b(b1_19to2_19),  .out_a(a2_19to2_20), .out_b(b2_19to3_19), .out_c(matrixC2_19));
processing_element pe2_20(.reset(effective_rst), .clk(clk),  .in_a(a2_19to2_20), .in_b(b1_20to2_20),  .out_a(a2_20to2_21), .out_b(b2_20to3_20), .out_c(matrixC2_20));
processing_element pe2_21(.reset(effective_rst), .clk(clk),  .in_a(a2_20to2_21), .in_b(b1_21to2_21),  .out_a(a2_21to2_22), .out_b(b2_21to3_21), .out_c(matrixC2_21));
processing_element pe2_22(.reset(effective_rst), .clk(clk),  .in_a(a2_21to2_22), .in_b(b1_22to2_22),  .out_a(a2_22to2_23), .out_b(b2_22to3_22), .out_c(matrixC2_22));
processing_element pe2_23(.reset(effective_rst), .clk(clk),  .in_a(a2_22to2_23), .in_b(b1_23to2_23),  .out_a(a2_23to2_24), .out_b(b2_23to3_23), .out_c(matrixC2_23));
processing_element pe2_24(.reset(effective_rst), .clk(clk),  .in_a(a2_23to2_24), .in_b(b1_24to2_24),  .out_a(a2_24to2_25), .out_b(b2_24to3_24), .out_c(matrixC2_24));
processing_element pe2_25(.reset(effective_rst), .clk(clk),  .in_a(a2_24to2_25), .in_b(b1_25to2_25),  .out_a(a2_25to2_26), .out_b(b2_25to3_25), .out_c(matrixC2_25));
processing_element pe2_26(.reset(effective_rst), .clk(clk),  .in_a(a2_25to2_26), .in_b(b1_26to2_26),  .out_a(a2_26to2_27), .out_b(b2_26to3_26), .out_c(matrixC2_26));
processing_element pe2_27(.reset(effective_rst), .clk(clk),  .in_a(a2_26to2_27), .in_b(b1_27to2_27),  .out_a(a2_27to2_28), .out_b(b2_27to3_27), .out_c(matrixC2_27));
processing_element pe2_28(.reset(effective_rst), .clk(clk),  .in_a(a2_27to2_28), .in_b(b1_28to2_28),  .out_a(a2_28to2_29), .out_b(b2_28to3_28), .out_c(matrixC2_28));
processing_element pe2_29(.reset(effective_rst), .clk(clk),  .in_a(a2_28to2_29), .in_b(b1_29to2_29),  .out_a(a2_29to2_30), .out_b(b2_29to3_29), .out_c(matrixC2_29));
processing_element pe2_30(.reset(effective_rst), .clk(clk),  .in_a(a2_29to2_30), .in_b(b1_30to2_30),  .out_a(a2_30to2_31), .out_b(b2_30to3_30), .out_c(matrixC2_30));
processing_element pe2_31(.reset(effective_rst), .clk(clk),  .in_a(a2_30to2_31), .in_b(b1_31to2_31),  .out_a(a2_31to2_32), .out_b(b2_31to3_31), .out_c(matrixC2_31));
processing_element pe3_1(.reset(effective_rst), .clk(clk),  .in_a(a3_0to3_1), .in_b(b2_1to3_1),  .out_a(a3_1to3_2), .out_b(b3_1to4_1), .out_c(matrixC3_1));
processing_element pe3_2(.reset(effective_rst), .clk(clk),  .in_a(a3_1to3_2), .in_b(b2_2to3_2),  .out_a(a3_2to3_3), .out_b(b3_2to4_2), .out_c(matrixC3_2));
processing_element pe3_3(.reset(effective_rst), .clk(clk),  .in_a(a3_2to3_3), .in_b(b2_3to3_3),  .out_a(a3_3to3_4), .out_b(b3_3to4_3), .out_c(matrixC3_3));
processing_element pe3_4(.reset(effective_rst), .clk(clk),  .in_a(a3_3to3_4), .in_b(b2_4to3_4),  .out_a(a3_4to3_5), .out_b(b3_4to4_4), .out_c(matrixC3_4));
processing_element pe3_5(.reset(effective_rst), .clk(clk),  .in_a(a3_4to3_5), .in_b(b2_5to3_5),  .out_a(a3_5to3_6), .out_b(b3_5to4_5), .out_c(matrixC3_5));
processing_element pe3_6(.reset(effective_rst), .clk(clk),  .in_a(a3_5to3_6), .in_b(b2_6to3_6),  .out_a(a3_6to3_7), .out_b(b3_6to4_6), .out_c(matrixC3_6));
processing_element pe3_7(.reset(effective_rst), .clk(clk),  .in_a(a3_6to3_7), .in_b(b2_7to3_7),  .out_a(a3_7to3_8), .out_b(b3_7to4_7), .out_c(matrixC3_7));
processing_element pe3_8(.reset(effective_rst), .clk(clk),  .in_a(a3_7to3_8), .in_b(b2_8to3_8),  .out_a(a3_8to3_9), .out_b(b3_8to4_8), .out_c(matrixC3_8));
processing_element pe3_9(.reset(effective_rst), .clk(clk),  .in_a(a3_8to3_9), .in_b(b2_9to3_9),  .out_a(a3_9to3_10), .out_b(b3_9to4_9), .out_c(matrixC3_9));
processing_element pe3_10(.reset(effective_rst), .clk(clk),  .in_a(a3_9to3_10), .in_b(b2_10to3_10),  .out_a(a3_10to3_11), .out_b(b3_10to4_10), .out_c(matrixC3_10));
processing_element pe3_11(.reset(effective_rst), .clk(clk),  .in_a(a3_10to3_11), .in_b(b2_11to3_11),  .out_a(a3_11to3_12), .out_b(b3_11to4_11), .out_c(matrixC3_11));
processing_element pe3_12(.reset(effective_rst), .clk(clk),  .in_a(a3_11to3_12), .in_b(b2_12to3_12),  .out_a(a3_12to3_13), .out_b(b3_12to4_12), .out_c(matrixC3_12));
processing_element pe3_13(.reset(effective_rst), .clk(clk),  .in_a(a3_12to3_13), .in_b(b2_13to3_13),  .out_a(a3_13to3_14), .out_b(b3_13to4_13), .out_c(matrixC3_13));
processing_element pe3_14(.reset(effective_rst), .clk(clk),  .in_a(a3_13to3_14), .in_b(b2_14to3_14),  .out_a(a3_14to3_15), .out_b(b3_14to4_14), .out_c(matrixC3_14));
processing_element pe3_15(.reset(effective_rst), .clk(clk),  .in_a(a3_14to3_15), .in_b(b2_15to3_15),  .out_a(a3_15to3_16), .out_b(b3_15to4_15), .out_c(matrixC3_15));
processing_element pe3_16(.reset(effective_rst), .clk(clk),  .in_a(a3_15to3_16), .in_b(b2_16to3_16),  .out_a(a3_16to3_17), .out_b(b3_16to4_16), .out_c(matrixC3_16));
processing_element pe3_17(.reset(effective_rst), .clk(clk),  .in_a(a3_16to3_17), .in_b(b2_17to3_17),  .out_a(a3_17to3_18), .out_b(b3_17to4_17), .out_c(matrixC3_17));
processing_element pe3_18(.reset(effective_rst), .clk(clk),  .in_a(a3_17to3_18), .in_b(b2_18to3_18),  .out_a(a3_18to3_19), .out_b(b3_18to4_18), .out_c(matrixC3_18));
processing_element pe3_19(.reset(effective_rst), .clk(clk),  .in_a(a3_18to3_19), .in_b(b2_19to3_19),  .out_a(a3_19to3_20), .out_b(b3_19to4_19), .out_c(matrixC3_19));
processing_element pe3_20(.reset(effective_rst), .clk(clk),  .in_a(a3_19to3_20), .in_b(b2_20to3_20),  .out_a(a3_20to3_21), .out_b(b3_20to4_20), .out_c(matrixC3_20));
processing_element pe3_21(.reset(effective_rst), .clk(clk),  .in_a(a3_20to3_21), .in_b(b2_21to3_21),  .out_a(a3_21to3_22), .out_b(b3_21to4_21), .out_c(matrixC3_21));
processing_element pe3_22(.reset(effective_rst), .clk(clk),  .in_a(a3_21to3_22), .in_b(b2_22to3_22),  .out_a(a3_22to3_23), .out_b(b3_22to4_22), .out_c(matrixC3_22));
processing_element pe3_23(.reset(effective_rst), .clk(clk),  .in_a(a3_22to3_23), .in_b(b2_23to3_23),  .out_a(a3_23to3_24), .out_b(b3_23to4_23), .out_c(matrixC3_23));
processing_element pe3_24(.reset(effective_rst), .clk(clk),  .in_a(a3_23to3_24), .in_b(b2_24to3_24),  .out_a(a3_24to3_25), .out_b(b3_24to4_24), .out_c(matrixC3_24));
processing_element pe3_25(.reset(effective_rst), .clk(clk),  .in_a(a3_24to3_25), .in_b(b2_25to3_25),  .out_a(a3_25to3_26), .out_b(b3_25to4_25), .out_c(matrixC3_25));
processing_element pe3_26(.reset(effective_rst), .clk(clk),  .in_a(a3_25to3_26), .in_b(b2_26to3_26),  .out_a(a3_26to3_27), .out_b(b3_26to4_26), .out_c(matrixC3_26));
processing_element pe3_27(.reset(effective_rst), .clk(clk),  .in_a(a3_26to3_27), .in_b(b2_27to3_27),  .out_a(a3_27to3_28), .out_b(b3_27to4_27), .out_c(matrixC3_27));
processing_element pe3_28(.reset(effective_rst), .clk(clk),  .in_a(a3_27to3_28), .in_b(b2_28to3_28),  .out_a(a3_28to3_29), .out_b(b3_28to4_28), .out_c(matrixC3_28));
processing_element pe3_29(.reset(effective_rst), .clk(clk),  .in_a(a3_28to3_29), .in_b(b2_29to3_29),  .out_a(a3_29to3_30), .out_b(b3_29to4_29), .out_c(matrixC3_29));
processing_element pe3_30(.reset(effective_rst), .clk(clk),  .in_a(a3_29to3_30), .in_b(b2_30to3_30),  .out_a(a3_30to3_31), .out_b(b3_30to4_30), .out_c(matrixC3_30));
processing_element pe3_31(.reset(effective_rst), .clk(clk),  .in_a(a3_30to3_31), .in_b(b2_31to3_31),  .out_a(a3_31to3_32), .out_b(b3_31to4_31), .out_c(matrixC3_31));
processing_element pe4_1(.reset(effective_rst), .clk(clk),  .in_a(a4_0to4_1), .in_b(b3_1to4_1),  .out_a(a4_1to4_2), .out_b(b4_1to5_1), .out_c(matrixC4_1));
processing_element pe4_2(.reset(effective_rst), .clk(clk),  .in_a(a4_1to4_2), .in_b(b3_2to4_2),  .out_a(a4_2to4_3), .out_b(b4_2to5_2), .out_c(matrixC4_2));
processing_element pe4_3(.reset(effective_rst), .clk(clk),  .in_a(a4_2to4_3), .in_b(b3_3to4_3),  .out_a(a4_3to4_4), .out_b(b4_3to5_3), .out_c(matrixC4_3));
processing_element pe4_4(.reset(effective_rst), .clk(clk),  .in_a(a4_3to4_4), .in_b(b3_4to4_4),  .out_a(a4_4to4_5), .out_b(b4_4to5_4), .out_c(matrixC4_4));
processing_element pe4_5(.reset(effective_rst), .clk(clk),  .in_a(a4_4to4_5), .in_b(b3_5to4_5),  .out_a(a4_5to4_6), .out_b(b4_5to5_5), .out_c(matrixC4_5));
processing_element pe4_6(.reset(effective_rst), .clk(clk),  .in_a(a4_5to4_6), .in_b(b3_6to4_6),  .out_a(a4_6to4_7), .out_b(b4_6to5_6), .out_c(matrixC4_6));
processing_element pe4_7(.reset(effective_rst), .clk(clk),  .in_a(a4_6to4_7), .in_b(b3_7to4_7),  .out_a(a4_7to4_8), .out_b(b4_7to5_7), .out_c(matrixC4_7));
processing_element pe4_8(.reset(effective_rst), .clk(clk),  .in_a(a4_7to4_8), .in_b(b3_8to4_8),  .out_a(a4_8to4_9), .out_b(b4_8to5_8), .out_c(matrixC4_8));
processing_element pe4_9(.reset(effective_rst), .clk(clk),  .in_a(a4_8to4_9), .in_b(b3_9to4_9),  .out_a(a4_9to4_10), .out_b(b4_9to5_9), .out_c(matrixC4_9));
processing_element pe4_10(.reset(effective_rst), .clk(clk),  .in_a(a4_9to4_10), .in_b(b3_10to4_10),  .out_a(a4_10to4_11), .out_b(b4_10to5_10), .out_c(matrixC4_10));
processing_element pe4_11(.reset(effective_rst), .clk(clk),  .in_a(a4_10to4_11), .in_b(b3_11to4_11),  .out_a(a4_11to4_12), .out_b(b4_11to5_11), .out_c(matrixC4_11));
processing_element pe4_12(.reset(effective_rst), .clk(clk),  .in_a(a4_11to4_12), .in_b(b3_12to4_12),  .out_a(a4_12to4_13), .out_b(b4_12to5_12), .out_c(matrixC4_12));
processing_element pe4_13(.reset(effective_rst), .clk(clk),  .in_a(a4_12to4_13), .in_b(b3_13to4_13),  .out_a(a4_13to4_14), .out_b(b4_13to5_13), .out_c(matrixC4_13));
processing_element pe4_14(.reset(effective_rst), .clk(clk),  .in_a(a4_13to4_14), .in_b(b3_14to4_14),  .out_a(a4_14to4_15), .out_b(b4_14to5_14), .out_c(matrixC4_14));
processing_element pe4_15(.reset(effective_rst), .clk(clk),  .in_a(a4_14to4_15), .in_b(b3_15to4_15),  .out_a(a4_15to4_16), .out_b(b4_15to5_15), .out_c(matrixC4_15));
processing_element pe4_16(.reset(effective_rst), .clk(clk),  .in_a(a4_15to4_16), .in_b(b3_16to4_16),  .out_a(a4_16to4_17), .out_b(b4_16to5_16), .out_c(matrixC4_16));
processing_element pe4_17(.reset(effective_rst), .clk(clk),  .in_a(a4_16to4_17), .in_b(b3_17to4_17),  .out_a(a4_17to4_18), .out_b(b4_17to5_17), .out_c(matrixC4_17));
processing_element pe4_18(.reset(effective_rst), .clk(clk),  .in_a(a4_17to4_18), .in_b(b3_18to4_18),  .out_a(a4_18to4_19), .out_b(b4_18to5_18), .out_c(matrixC4_18));
processing_element pe4_19(.reset(effective_rst), .clk(clk),  .in_a(a4_18to4_19), .in_b(b3_19to4_19),  .out_a(a4_19to4_20), .out_b(b4_19to5_19), .out_c(matrixC4_19));
processing_element pe4_20(.reset(effective_rst), .clk(clk),  .in_a(a4_19to4_20), .in_b(b3_20to4_20),  .out_a(a4_20to4_21), .out_b(b4_20to5_20), .out_c(matrixC4_20));
processing_element pe4_21(.reset(effective_rst), .clk(clk),  .in_a(a4_20to4_21), .in_b(b3_21to4_21),  .out_a(a4_21to4_22), .out_b(b4_21to5_21), .out_c(matrixC4_21));
processing_element pe4_22(.reset(effective_rst), .clk(clk),  .in_a(a4_21to4_22), .in_b(b3_22to4_22),  .out_a(a4_22to4_23), .out_b(b4_22to5_22), .out_c(matrixC4_22));
processing_element pe4_23(.reset(effective_rst), .clk(clk),  .in_a(a4_22to4_23), .in_b(b3_23to4_23),  .out_a(a4_23to4_24), .out_b(b4_23to5_23), .out_c(matrixC4_23));
processing_element pe4_24(.reset(effective_rst), .clk(clk),  .in_a(a4_23to4_24), .in_b(b3_24to4_24),  .out_a(a4_24to4_25), .out_b(b4_24to5_24), .out_c(matrixC4_24));
processing_element pe4_25(.reset(effective_rst), .clk(clk),  .in_a(a4_24to4_25), .in_b(b3_25to4_25),  .out_a(a4_25to4_26), .out_b(b4_25to5_25), .out_c(matrixC4_25));
processing_element pe4_26(.reset(effective_rst), .clk(clk),  .in_a(a4_25to4_26), .in_b(b3_26to4_26),  .out_a(a4_26to4_27), .out_b(b4_26to5_26), .out_c(matrixC4_26));
processing_element pe4_27(.reset(effective_rst), .clk(clk),  .in_a(a4_26to4_27), .in_b(b3_27to4_27),  .out_a(a4_27to4_28), .out_b(b4_27to5_27), .out_c(matrixC4_27));
processing_element pe4_28(.reset(effective_rst), .clk(clk),  .in_a(a4_27to4_28), .in_b(b3_28to4_28),  .out_a(a4_28to4_29), .out_b(b4_28to5_28), .out_c(matrixC4_28));
processing_element pe4_29(.reset(effective_rst), .clk(clk),  .in_a(a4_28to4_29), .in_b(b3_29to4_29),  .out_a(a4_29to4_30), .out_b(b4_29to5_29), .out_c(matrixC4_29));
processing_element pe4_30(.reset(effective_rst), .clk(clk),  .in_a(a4_29to4_30), .in_b(b3_30to4_30),  .out_a(a4_30to4_31), .out_b(b4_30to5_30), .out_c(matrixC4_30));
processing_element pe4_31(.reset(effective_rst), .clk(clk),  .in_a(a4_30to4_31), .in_b(b3_31to4_31),  .out_a(a4_31to4_32), .out_b(b4_31to5_31), .out_c(matrixC4_31));
processing_element pe5_1(.reset(effective_rst), .clk(clk),  .in_a(a5_0to5_1), .in_b(b4_1to5_1),  .out_a(a5_1to5_2), .out_b(b5_1to6_1), .out_c(matrixC5_1));
processing_element pe5_2(.reset(effective_rst), .clk(clk),  .in_a(a5_1to5_2), .in_b(b4_2to5_2),  .out_a(a5_2to5_3), .out_b(b5_2to6_2), .out_c(matrixC5_2));
processing_element pe5_3(.reset(effective_rst), .clk(clk),  .in_a(a5_2to5_3), .in_b(b4_3to5_3),  .out_a(a5_3to5_4), .out_b(b5_3to6_3), .out_c(matrixC5_3));
processing_element pe5_4(.reset(effective_rst), .clk(clk),  .in_a(a5_3to5_4), .in_b(b4_4to5_4),  .out_a(a5_4to5_5), .out_b(b5_4to6_4), .out_c(matrixC5_4));
processing_element pe5_5(.reset(effective_rst), .clk(clk),  .in_a(a5_4to5_5), .in_b(b4_5to5_5),  .out_a(a5_5to5_6), .out_b(b5_5to6_5), .out_c(matrixC5_5));
processing_element pe5_6(.reset(effective_rst), .clk(clk),  .in_a(a5_5to5_6), .in_b(b4_6to5_6),  .out_a(a5_6to5_7), .out_b(b5_6to6_6), .out_c(matrixC5_6));
processing_element pe5_7(.reset(effective_rst), .clk(clk),  .in_a(a5_6to5_7), .in_b(b4_7to5_7),  .out_a(a5_7to5_8), .out_b(b5_7to6_7), .out_c(matrixC5_7));
processing_element pe5_8(.reset(effective_rst), .clk(clk),  .in_a(a5_7to5_8), .in_b(b4_8to5_8),  .out_a(a5_8to5_9), .out_b(b5_8to6_8), .out_c(matrixC5_8));
processing_element pe5_9(.reset(effective_rst), .clk(clk),  .in_a(a5_8to5_9), .in_b(b4_9to5_9),  .out_a(a5_9to5_10), .out_b(b5_9to6_9), .out_c(matrixC5_9));
processing_element pe5_10(.reset(effective_rst), .clk(clk),  .in_a(a5_9to5_10), .in_b(b4_10to5_10),  .out_a(a5_10to5_11), .out_b(b5_10to6_10), .out_c(matrixC5_10));
processing_element pe5_11(.reset(effective_rst), .clk(clk),  .in_a(a5_10to5_11), .in_b(b4_11to5_11),  .out_a(a5_11to5_12), .out_b(b5_11to6_11), .out_c(matrixC5_11));
processing_element pe5_12(.reset(effective_rst), .clk(clk),  .in_a(a5_11to5_12), .in_b(b4_12to5_12),  .out_a(a5_12to5_13), .out_b(b5_12to6_12), .out_c(matrixC5_12));
processing_element pe5_13(.reset(effective_rst), .clk(clk),  .in_a(a5_12to5_13), .in_b(b4_13to5_13),  .out_a(a5_13to5_14), .out_b(b5_13to6_13), .out_c(matrixC5_13));
processing_element pe5_14(.reset(effective_rst), .clk(clk),  .in_a(a5_13to5_14), .in_b(b4_14to5_14),  .out_a(a5_14to5_15), .out_b(b5_14to6_14), .out_c(matrixC5_14));
processing_element pe5_15(.reset(effective_rst), .clk(clk),  .in_a(a5_14to5_15), .in_b(b4_15to5_15),  .out_a(a5_15to5_16), .out_b(b5_15to6_15), .out_c(matrixC5_15));
processing_element pe5_16(.reset(effective_rst), .clk(clk),  .in_a(a5_15to5_16), .in_b(b4_16to5_16),  .out_a(a5_16to5_17), .out_b(b5_16to6_16), .out_c(matrixC5_16));
processing_element pe5_17(.reset(effective_rst), .clk(clk),  .in_a(a5_16to5_17), .in_b(b4_17to5_17),  .out_a(a5_17to5_18), .out_b(b5_17to6_17), .out_c(matrixC5_17));
processing_element pe5_18(.reset(effective_rst), .clk(clk),  .in_a(a5_17to5_18), .in_b(b4_18to5_18),  .out_a(a5_18to5_19), .out_b(b5_18to6_18), .out_c(matrixC5_18));
processing_element pe5_19(.reset(effective_rst), .clk(clk),  .in_a(a5_18to5_19), .in_b(b4_19to5_19),  .out_a(a5_19to5_20), .out_b(b5_19to6_19), .out_c(matrixC5_19));
processing_element pe5_20(.reset(effective_rst), .clk(clk),  .in_a(a5_19to5_20), .in_b(b4_20to5_20),  .out_a(a5_20to5_21), .out_b(b5_20to6_20), .out_c(matrixC5_20));
processing_element pe5_21(.reset(effective_rst), .clk(clk),  .in_a(a5_20to5_21), .in_b(b4_21to5_21),  .out_a(a5_21to5_22), .out_b(b5_21to6_21), .out_c(matrixC5_21));
processing_element pe5_22(.reset(effective_rst), .clk(clk),  .in_a(a5_21to5_22), .in_b(b4_22to5_22),  .out_a(a5_22to5_23), .out_b(b5_22to6_22), .out_c(matrixC5_22));
processing_element pe5_23(.reset(effective_rst), .clk(clk),  .in_a(a5_22to5_23), .in_b(b4_23to5_23),  .out_a(a5_23to5_24), .out_b(b5_23to6_23), .out_c(matrixC5_23));
processing_element pe5_24(.reset(effective_rst), .clk(clk),  .in_a(a5_23to5_24), .in_b(b4_24to5_24),  .out_a(a5_24to5_25), .out_b(b5_24to6_24), .out_c(matrixC5_24));
processing_element pe5_25(.reset(effective_rst), .clk(clk),  .in_a(a5_24to5_25), .in_b(b4_25to5_25),  .out_a(a5_25to5_26), .out_b(b5_25to6_25), .out_c(matrixC5_25));
processing_element pe5_26(.reset(effective_rst), .clk(clk),  .in_a(a5_25to5_26), .in_b(b4_26to5_26),  .out_a(a5_26to5_27), .out_b(b5_26to6_26), .out_c(matrixC5_26));
processing_element pe5_27(.reset(effective_rst), .clk(clk),  .in_a(a5_26to5_27), .in_b(b4_27to5_27),  .out_a(a5_27to5_28), .out_b(b5_27to6_27), .out_c(matrixC5_27));
processing_element pe5_28(.reset(effective_rst), .clk(clk),  .in_a(a5_27to5_28), .in_b(b4_28to5_28),  .out_a(a5_28to5_29), .out_b(b5_28to6_28), .out_c(matrixC5_28));
processing_element pe5_29(.reset(effective_rst), .clk(clk),  .in_a(a5_28to5_29), .in_b(b4_29to5_29),  .out_a(a5_29to5_30), .out_b(b5_29to6_29), .out_c(matrixC5_29));
processing_element pe5_30(.reset(effective_rst), .clk(clk),  .in_a(a5_29to5_30), .in_b(b4_30to5_30),  .out_a(a5_30to5_31), .out_b(b5_30to6_30), .out_c(matrixC5_30));
processing_element pe5_31(.reset(effective_rst), .clk(clk),  .in_a(a5_30to5_31), .in_b(b4_31to5_31),  .out_a(a5_31to5_32), .out_b(b5_31to6_31), .out_c(matrixC5_31));
processing_element pe6_1(.reset(effective_rst), .clk(clk),  .in_a(a6_0to6_1), .in_b(b5_1to6_1),  .out_a(a6_1to6_2), .out_b(b6_1to7_1), .out_c(matrixC6_1));
processing_element pe6_2(.reset(effective_rst), .clk(clk),  .in_a(a6_1to6_2), .in_b(b5_2to6_2),  .out_a(a6_2to6_3), .out_b(b6_2to7_2), .out_c(matrixC6_2));
processing_element pe6_3(.reset(effective_rst), .clk(clk),  .in_a(a6_2to6_3), .in_b(b5_3to6_3),  .out_a(a6_3to6_4), .out_b(b6_3to7_3), .out_c(matrixC6_3));
processing_element pe6_4(.reset(effective_rst), .clk(clk),  .in_a(a6_3to6_4), .in_b(b5_4to6_4),  .out_a(a6_4to6_5), .out_b(b6_4to7_4), .out_c(matrixC6_4));
processing_element pe6_5(.reset(effective_rst), .clk(clk),  .in_a(a6_4to6_5), .in_b(b5_5to6_5),  .out_a(a6_5to6_6), .out_b(b6_5to7_5), .out_c(matrixC6_5));
processing_element pe6_6(.reset(effective_rst), .clk(clk),  .in_a(a6_5to6_6), .in_b(b5_6to6_6),  .out_a(a6_6to6_7), .out_b(b6_6to7_6), .out_c(matrixC6_6));
processing_element pe6_7(.reset(effective_rst), .clk(clk),  .in_a(a6_6to6_7), .in_b(b5_7to6_7),  .out_a(a6_7to6_8), .out_b(b6_7to7_7), .out_c(matrixC6_7));
processing_element pe6_8(.reset(effective_rst), .clk(clk),  .in_a(a6_7to6_8), .in_b(b5_8to6_8),  .out_a(a6_8to6_9), .out_b(b6_8to7_8), .out_c(matrixC6_8));
processing_element pe6_9(.reset(effective_rst), .clk(clk),  .in_a(a6_8to6_9), .in_b(b5_9to6_9),  .out_a(a6_9to6_10), .out_b(b6_9to7_9), .out_c(matrixC6_9));
processing_element pe6_10(.reset(effective_rst), .clk(clk),  .in_a(a6_9to6_10), .in_b(b5_10to6_10),  .out_a(a6_10to6_11), .out_b(b6_10to7_10), .out_c(matrixC6_10));
processing_element pe6_11(.reset(effective_rst), .clk(clk),  .in_a(a6_10to6_11), .in_b(b5_11to6_11),  .out_a(a6_11to6_12), .out_b(b6_11to7_11), .out_c(matrixC6_11));
processing_element pe6_12(.reset(effective_rst), .clk(clk),  .in_a(a6_11to6_12), .in_b(b5_12to6_12),  .out_a(a6_12to6_13), .out_b(b6_12to7_12), .out_c(matrixC6_12));
processing_element pe6_13(.reset(effective_rst), .clk(clk),  .in_a(a6_12to6_13), .in_b(b5_13to6_13),  .out_a(a6_13to6_14), .out_b(b6_13to7_13), .out_c(matrixC6_13));
processing_element pe6_14(.reset(effective_rst), .clk(clk),  .in_a(a6_13to6_14), .in_b(b5_14to6_14),  .out_a(a6_14to6_15), .out_b(b6_14to7_14), .out_c(matrixC6_14));
processing_element pe6_15(.reset(effective_rst), .clk(clk),  .in_a(a6_14to6_15), .in_b(b5_15to6_15),  .out_a(a6_15to6_16), .out_b(b6_15to7_15), .out_c(matrixC6_15));
processing_element pe6_16(.reset(effective_rst), .clk(clk),  .in_a(a6_15to6_16), .in_b(b5_16to6_16),  .out_a(a6_16to6_17), .out_b(b6_16to7_16), .out_c(matrixC6_16));
processing_element pe6_17(.reset(effective_rst), .clk(clk),  .in_a(a6_16to6_17), .in_b(b5_17to6_17),  .out_a(a6_17to6_18), .out_b(b6_17to7_17), .out_c(matrixC6_17));
processing_element pe6_18(.reset(effective_rst), .clk(clk),  .in_a(a6_17to6_18), .in_b(b5_18to6_18),  .out_a(a6_18to6_19), .out_b(b6_18to7_18), .out_c(matrixC6_18));
processing_element pe6_19(.reset(effective_rst), .clk(clk),  .in_a(a6_18to6_19), .in_b(b5_19to6_19),  .out_a(a6_19to6_20), .out_b(b6_19to7_19), .out_c(matrixC6_19));
processing_element pe6_20(.reset(effective_rst), .clk(clk),  .in_a(a6_19to6_20), .in_b(b5_20to6_20),  .out_a(a6_20to6_21), .out_b(b6_20to7_20), .out_c(matrixC6_20));
processing_element pe6_21(.reset(effective_rst), .clk(clk),  .in_a(a6_20to6_21), .in_b(b5_21to6_21),  .out_a(a6_21to6_22), .out_b(b6_21to7_21), .out_c(matrixC6_21));
processing_element pe6_22(.reset(effective_rst), .clk(clk),  .in_a(a6_21to6_22), .in_b(b5_22to6_22),  .out_a(a6_22to6_23), .out_b(b6_22to7_22), .out_c(matrixC6_22));
processing_element pe6_23(.reset(effective_rst), .clk(clk),  .in_a(a6_22to6_23), .in_b(b5_23to6_23),  .out_a(a6_23to6_24), .out_b(b6_23to7_23), .out_c(matrixC6_23));
processing_element pe6_24(.reset(effective_rst), .clk(clk),  .in_a(a6_23to6_24), .in_b(b5_24to6_24),  .out_a(a6_24to6_25), .out_b(b6_24to7_24), .out_c(matrixC6_24));
processing_element pe6_25(.reset(effective_rst), .clk(clk),  .in_a(a6_24to6_25), .in_b(b5_25to6_25),  .out_a(a6_25to6_26), .out_b(b6_25to7_25), .out_c(matrixC6_25));
processing_element pe6_26(.reset(effective_rst), .clk(clk),  .in_a(a6_25to6_26), .in_b(b5_26to6_26),  .out_a(a6_26to6_27), .out_b(b6_26to7_26), .out_c(matrixC6_26));
processing_element pe6_27(.reset(effective_rst), .clk(clk),  .in_a(a6_26to6_27), .in_b(b5_27to6_27),  .out_a(a6_27to6_28), .out_b(b6_27to7_27), .out_c(matrixC6_27));
processing_element pe6_28(.reset(effective_rst), .clk(clk),  .in_a(a6_27to6_28), .in_b(b5_28to6_28),  .out_a(a6_28to6_29), .out_b(b6_28to7_28), .out_c(matrixC6_28));
processing_element pe6_29(.reset(effective_rst), .clk(clk),  .in_a(a6_28to6_29), .in_b(b5_29to6_29),  .out_a(a6_29to6_30), .out_b(b6_29to7_29), .out_c(matrixC6_29));
processing_element pe6_30(.reset(effective_rst), .clk(clk),  .in_a(a6_29to6_30), .in_b(b5_30to6_30),  .out_a(a6_30to6_31), .out_b(b6_30to7_30), .out_c(matrixC6_30));
processing_element pe6_31(.reset(effective_rst), .clk(clk),  .in_a(a6_30to6_31), .in_b(b5_31to6_31),  .out_a(a6_31to6_32), .out_b(b6_31to7_31), .out_c(matrixC6_31));
processing_element pe7_1(.reset(effective_rst), .clk(clk),  .in_a(a7_0to7_1), .in_b(b6_1to7_1),  .out_a(a7_1to7_2), .out_b(b7_1to8_1), .out_c(matrixC7_1));
processing_element pe7_2(.reset(effective_rst), .clk(clk),  .in_a(a7_1to7_2), .in_b(b6_2to7_2),  .out_a(a7_2to7_3), .out_b(b7_2to8_2), .out_c(matrixC7_2));
processing_element pe7_3(.reset(effective_rst), .clk(clk),  .in_a(a7_2to7_3), .in_b(b6_3to7_3),  .out_a(a7_3to7_4), .out_b(b7_3to8_3), .out_c(matrixC7_3));
processing_element pe7_4(.reset(effective_rst), .clk(clk),  .in_a(a7_3to7_4), .in_b(b6_4to7_4),  .out_a(a7_4to7_5), .out_b(b7_4to8_4), .out_c(matrixC7_4));
processing_element pe7_5(.reset(effective_rst), .clk(clk),  .in_a(a7_4to7_5), .in_b(b6_5to7_5),  .out_a(a7_5to7_6), .out_b(b7_5to8_5), .out_c(matrixC7_5));
processing_element pe7_6(.reset(effective_rst), .clk(clk),  .in_a(a7_5to7_6), .in_b(b6_6to7_6),  .out_a(a7_6to7_7), .out_b(b7_6to8_6), .out_c(matrixC7_6));
processing_element pe7_7(.reset(effective_rst), .clk(clk),  .in_a(a7_6to7_7), .in_b(b6_7to7_7),  .out_a(a7_7to7_8), .out_b(b7_7to8_7), .out_c(matrixC7_7));
processing_element pe7_8(.reset(effective_rst), .clk(clk),  .in_a(a7_7to7_8), .in_b(b6_8to7_8),  .out_a(a7_8to7_9), .out_b(b7_8to8_8), .out_c(matrixC7_8));
processing_element pe7_9(.reset(effective_rst), .clk(clk),  .in_a(a7_8to7_9), .in_b(b6_9to7_9),  .out_a(a7_9to7_10), .out_b(b7_9to8_9), .out_c(matrixC7_9));
processing_element pe7_10(.reset(effective_rst), .clk(clk),  .in_a(a7_9to7_10), .in_b(b6_10to7_10),  .out_a(a7_10to7_11), .out_b(b7_10to8_10), .out_c(matrixC7_10));
processing_element pe7_11(.reset(effective_rst), .clk(clk),  .in_a(a7_10to7_11), .in_b(b6_11to7_11),  .out_a(a7_11to7_12), .out_b(b7_11to8_11), .out_c(matrixC7_11));
processing_element pe7_12(.reset(effective_rst), .clk(clk),  .in_a(a7_11to7_12), .in_b(b6_12to7_12),  .out_a(a7_12to7_13), .out_b(b7_12to8_12), .out_c(matrixC7_12));
processing_element pe7_13(.reset(effective_rst), .clk(clk),  .in_a(a7_12to7_13), .in_b(b6_13to7_13),  .out_a(a7_13to7_14), .out_b(b7_13to8_13), .out_c(matrixC7_13));
processing_element pe7_14(.reset(effective_rst), .clk(clk),  .in_a(a7_13to7_14), .in_b(b6_14to7_14),  .out_a(a7_14to7_15), .out_b(b7_14to8_14), .out_c(matrixC7_14));
processing_element pe7_15(.reset(effective_rst), .clk(clk),  .in_a(a7_14to7_15), .in_b(b6_15to7_15),  .out_a(a7_15to7_16), .out_b(b7_15to8_15), .out_c(matrixC7_15));
processing_element pe7_16(.reset(effective_rst), .clk(clk),  .in_a(a7_15to7_16), .in_b(b6_16to7_16),  .out_a(a7_16to7_17), .out_b(b7_16to8_16), .out_c(matrixC7_16));
processing_element pe7_17(.reset(effective_rst), .clk(clk),  .in_a(a7_16to7_17), .in_b(b6_17to7_17),  .out_a(a7_17to7_18), .out_b(b7_17to8_17), .out_c(matrixC7_17));
processing_element pe7_18(.reset(effective_rst), .clk(clk),  .in_a(a7_17to7_18), .in_b(b6_18to7_18),  .out_a(a7_18to7_19), .out_b(b7_18to8_18), .out_c(matrixC7_18));
processing_element pe7_19(.reset(effective_rst), .clk(clk),  .in_a(a7_18to7_19), .in_b(b6_19to7_19),  .out_a(a7_19to7_20), .out_b(b7_19to8_19), .out_c(matrixC7_19));
processing_element pe7_20(.reset(effective_rst), .clk(clk),  .in_a(a7_19to7_20), .in_b(b6_20to7_20),  .out_a(a7_20to7_21), .out_b(b7_20to8_20), .out_c(matrixC7_20));
processing_element pe7_21(.reset(effective_rst), .clk(clk),  .in_a(a7_20to7_21), .in_b(b6_21to7_21),  .out_a(a7_21to7_22), .out_b(b7_21to8_21), .out_c(matrixC7_21));
processing_element pe7_22(.reset(effective_rst), .clk(clk),  .in_a(a7_21to7_22), .in_b(b6_22to7_22),  .out_a(a7_22to7_23), .out_b(b7_22to8_22), .out_c(matrixC7_22));
processing_element pe7_23(.reset(effective_rst), .clk(clk),  .in_a(a7_22to7_23), .in_b(b6_23to7_23),  .out_a(a7_23to7_24), .out_b(b7_23to8_23), .out_c(matrixC7_23));
processing_element pe7_24(.reset(effective_rst), .clk(clk),  .in_a(a7_23to7_24), .in_b(b6_24to7_24),  .out_a(a7_24to7_25), .out_b(b7_24to8_24), .out_c(matrixC7_24));
processing_element pe7_25(.reset(effective_rst), .clk(clk),  .in_a(a7_24to7_25), .in_b(b6_25to7_25),  .out_a(a7_25to7_26), .out_b(b7_25to8_25), .out_c(matrixC7_25));
processing_element pe7_26(.reset(effective_rst), .clk(clk),  .in_a(a7_25to7_26), .in_b(b6_26to7_26),  .out_a(a7_26to7_27), .out_b(b7_26to8_26), .out_c(matrixC7_26));
processing_element pe7_27(.reset(effective_rst), .clk(clk),  .in_a(a7_26to7_27), .in_b(b6_27to7_27),  .out_a(a7_27to7_28), .out_b(b7_27to8_27), .out_c(matrixC7_27));
processing_element pe7_28(.reset(effective_rst), .clk(clk),  .in_a(a7_27to7_28), .in_b(b6_28to7_28),  .out_a(a7_28to7_29), .out_b(b7_28to8_28), .out_c(matrixC7_28));
processing_element pe7_29(.reset(effective_rst), .clk(clk),  .in_a(a7_28to7_29), .in_b(b6_29to7_29),  .out_a(a7_29to7_30), .out_b(b7_29to8_29), .out_c(matrixC7_29));
processing_element pe7_30(.reset(effective_rst), .clk(clk),  .in_a(a7_29to7_30), .in_b(b6_30to7_30),  .out_a(a7_30to7_31), .out_b(b7_30to8_30), .out_c(matrixC7_30));
processing_element pe7_31(.reset(effective_rst), .clk(clk),  .in_a(a7_30to7_31), .in_b(b6_31to7_31),  .out_a(a7_31to7_32), .out_b(b7_31to8_31), .out_c(matrixC7_31));
processing_element pe8_1(.reset(effective_rst), .clk(clk),  .in_a(a8_0to8_1), .in_b(b7_1to8_1),  .out_a(a8_1to8_2), .out_b(b8_1to9_1), .out_c(matrixC8_1));
processing_element pe8_2(.reset(effective_rst), .clk(clk),  .in_a(a8_1to8_2), .in_b(b7_2to8_2),  .out_a(a8_2to8_3), .out_b(b8_2to9_2), .out_c(matrixC8_2));
processing_element pe8_3(.reset(effective_rst), .clk(clk),  .in_a(a8_2to8_3), .in_b(b7_3to8_3),  .out_a(a8_3to8_4), .out_b(b8_3to9_3), .out_c(matrixC8_3));
processing_element pe8_4(.reset(effective_rst), .clk(clk),  .in_a(a8_3to8_4), .in_b(b7_4to8_4),  .out_a(a8_4to8_5), .out_b(b8_4to9_4), .out_c(matrixC8_4));
processing_element pe8_5(.reset(effective_rst), .clk(clk),  .in_a(a8_4to8_5), .in_b(b7_5to8_5),  .out_a(a8_5to8_6), .out_b(b8_5to9_5), .out_c(matrixC8_5));
processing_element pe8_6(.reset(effective_rst), .clk(clk),  .in_a(a8_5to8_6), .in_b(b7_6to8_6),  .out_a(a8_6to8_7), .out_b(b8_6to9_6), .out_c(matrixC8_6));
processing_element pe8_7(.reset(effective_rst), .clk(clk),  .in_a(a8_6to8_7), .in_b(b7_7to8_7),  .out_a(a8_7to8_8), .out_b(b8_7to9_7), .out_c(matrixC8_7));
processing_element pe8_8(.reset(effective_rst), .clk(clk),  .in_a(a8_7to8_8), .in_b(b7_8to8_8),  .out_a(a8_8to8_9), .out_b(b8_8to9_8), .out_c(matrixC8_8));
processing_element pe8_9(.reset(effective_rst), .clk(clk),  .in_a(a8_8to8_9), .in_b(b7_9to8_9),  .out_a(a8_9to8_10), .out_b(b8_9to9_9), .out_c(matrixC8_9));
processing_element pe8_10(.reset(effective_rst), .clk(clk),  .in_a(a8_9to8_10), .in_b(b7_10to8_10),  .out_a(a8_10to8_11), .out_b(b8_10to9_10), .out_c(matrixC8_10));
processing_element pe8_11(.reset(effective_rst), .clk(clk),  .in_a(a8_10to8_11), .in_b(b7_11to8_11),  .out_a(a8_11to8_12), .out_b(b8_11to9_11), .out_c(matrixC8_11));
processing_element pe8_12(.reset(effective_rst), .clk(clk),  .in_a(a8_11to8_12), .in_b(b7_12to8_12),  .out_a(a8_12to8_13), .out_b(b8_12to9_12), .out_c(matrixC8_12));
processing_element pe8_13(.reset(effective_rst), .clk(clk),  .in_a(a8_12to8_13), .in_b(b7_13to8_13),  .out_a(a8_13to8_14), .out_b(b8_13to9_13), .out_c(matrixC8_13));
processing_element pe8_14(.reset(effective_rst), .clk(clk),  .in_a(a8_13to8_14), .in_b(b7_14to8_14),  .out_a(a8_14to8_15), .out_b(b8_14to9_14), .out_c(matrixC8_14));
processing_element pe8_15(.reset(effective_rst), .clk(clk),  .in_a(a8_14to8_15), .in_b(b7_15to8_15),  .out_a(a8_15to8_16), .out_b(b8_15to9_15), .out_c(matrixC8_15));
processing_element pe8_16(.reset(effective_rst), .clk(clk),  .in_a(a8_15to8_16), .in_b(b7_16to8_16),  .out_a(a8_16to8_17), .out_b(b8_16to9_16), .out_c(matrixC8_16));
processing_element pe8_17(.reset(effective_rst), .clk(clk),  .in_a(a8_16to8_17), .in_b(b7_17to8_17),  .out_a(a8_17to8_18), .out_b(b8_17to9_17), .out_c(matrixC8_17));
processing_element pe8_18(.reset(effective_rst), .clk(clk),  .in_a(a8_17to8_18), .in_b(b7_18to8_18),  .out_a(a8_18to8_19), .out_b(b8_18to9_18), .out_c(matrixC8_18));
processing_element pe8_19(.reset(effective_rst), .clk(clk),  .in_a(a8_18to8_19), .in_b(b7_19to8_19),  .out_a(a8_19to8_20), .out_b(b8_19to9_19), .out_c(matrixC8_19));
processing_element pe8_20(.reset(effective_rst), .clk(clk),  .in_a(a8_19to8_20), .in_b(b7_20to8_20),  .out_a(a8_20to8_21), .out_b(b8_20to9_20), .out_c(matrixC8_20));
processing_element pe8_21(.reset(effective_rst), .clk(clk),  .in_a(a8_20to8_21), .in_b(b7_21to8_21),  .out_a(a8_21to8_22), .out_b(b8_21to9_21), .out_c(matrixC8_21));
processing_element pe8_22(.reset(effective_rst), .clk(clk),  .in_a(a8_21to8_22), .in_b(b7_22to8_22),  .out_a(a8_22to8_23), .out_b(b8_22to9_22), .out_c(matrixC8_22));
processing_element pe8_23(.reset(effective_rst), .clk(clk),  .in_a(a8_22to8_23), .in_b(b7_23to8_23),  .out_a(a8_23to8_24), .out_b(b8_23to9_23), .out_c(matrixC8_23));
processing_element pe8_24(.reset(effective_rst), .clk(clk),  .in_a(a8_23to8_24), .in_b(b7_24to8_24),  .out_a(a8_24to8_25), .out_b(b8_24to9_24), .out_c(matrixC8_24));
processing_element pe8_25(.reset(effective_rst), .clk(clk),  .in_a(a8_24to8_25), .in_b(b7_25to8_25),  .out_a(a8_25to8_26), .out_b(b8_25to9_25), .out_c(matrixC8_25));
processing_element pe8_26(.reset(effective_rst), .clk(clk),  .in_a(a8_25to8_26), .in_b(b7_26to8_26),  .out_a(a8_26to8_27), .out_b(b8_26to9_26), .out_c(matrixC8_26));
processing_element pe8_27(.reset(effective_rst), .clk(clk),  .in_a(a8_26to8_27), .in_b(b7_27to8_27),  .out_a(a8_27to8_28), .out_b(b8_27to9_27), .out_c(matrixC8_27));
processing_element pe8_28(.reset(effective_rst), .clk(clk),  .in_a(a8_27to8_28), .in_b(b7_28to8_28),  .out_a(a8_28to8_29), .out_b(b8_28to9_28), .out_c(matrixC8_28));
processing_element pe8_29(.reset(effective_rst), .clk(clk),  .in_a(a8_28to8_29), .in_b(b7_29to8_29),  .out_a(a8_29to8_30), .out_b(b8_29to9_29), .out_c(matrixC8_29));
processing_element pe8_30(.reset(effective_rst), .clk(clk),  .in_a(a8_29to8_30), .in_b(b7_30to8_30),  .out_a(a8_30to8_31), .out_b(b8_30to9_30), .out_c(matrixC8_30));
processing_element pe8_31(.reset(effective_rst), .clk(clk),  .in_a(a8_30to8_31), .in_b(b7_31to8_31),  .out_a(a8_31to8_32), .out_b(b8_31to9_31), .out_c(matrixC8_31));
processing_element pe9_1(.reset(effective_rst), .clk(clk),  .in_a(a9_0to9_1), .in_b(b8_1to9_1),  .out_a(a9_1to9_2), .out_b(b9_1to10_1), .out_c(matrixC9_1));
processing_element pe9_2(.reset(effective_rst), .clk(clk),  .in_a(a9_1to9_2), .in_b(b8_2to9_2),  .out_a(a9_2to9_3), .out_b(b9_2to10_2), .out_c(matrixC9_2));
processing_element pe9_3(.reset(effective_rst), .clk(clk),  .in_a(a9_2to9_3), .in_b(b8_3to9_3),  .out_a(a9_3to9_4), .out_b(b9_3to10_3), .out_c(matrixC9_3));
processing_element pe9_4(.reset(effective_rst), .clk(clk),  .in_a(a9_3to9_4), .in_b(b8_4to9_4),  .out_a(a9_4to9_5), .out_b(b9_4to10_4), .out_c(matrixC9_4));
processing_element pe9_5(.reset(effective_rst), .clk(clk),  .in_a(a9_4to9_5), .in_b(b8_5to9_5),  .out_a(a9_5to9_6), .out_b(b9_5to10_5), .out_c(matrixC9_5));
processing_element pe9_6(.reset(effective_rst), .clk(clk),  .in_a(a9_5to9_6), .in_b(b8_6to9_6),  .out_a(a9_6to9_7), .out_b(b9_6to10_6), .out_c(matrixC9_6));
processing_element pe9_7(.reset(effective_rst), .clk(clk),  .in_a(a9_6to9_7), .in_b(b8_7to9_7),  .out_a(a9_7to9_8), .out_b(b9_7to10_7), .out_c(matrixC9_7));
processing_element pe9_8(.reset(effective_rst), .clk(clk),  .in_a(a9_7to9_8), .in_b(b8_8to9_8),  .out_a(a9_8to9_9), .out_b(b9_8to10_8), .out_c(matrixC9_8));
processing_element pe9_9(.reset(effective_rst), .clk(clk),  .in_a(a9_8to9_9), .in_b(b8_9to9_9),  .out_a(a9_9to9_10), .out_b(b9_9to10_9), .out_c(matrixC9_9));
processing_element pe9_10(.reset(effective_rst), .clk(clk),  .in_a(a9_9to9_10), .in_b(b8_10to9_10),  .out_a(a9_10to9_11), .out_b(b9_10to10_10), .out_c(matrixC9_10));
processing_element pe9_11(.reset(effective_rst), .clk(clk),  .in_a(a9_10to9_11), .in_b(b8_11to9_11),  .out_a(a9_11to9_12), .out_b(b9_11to10_11), .out_c(matrixC9_11));
processing_element pe9_12(.reset(effective_rst), .clk(clk),  .in_a(a9_11to9_12), .in_b(b8_12to9_12),  .out_a(a9_12to9_13), .out_b(b9_12to10_12), .out_c(matrixC9_12));
processing_element pe9_13(.reset(effective_rst), .clk(clk),  .in_a(a9_12to9_13), .in_b(b8_13to9_13),  .out_a(a9_13to9_14), .out_b(b9_13to10_13), .out_c(matrixC9_13));
processing_element pe9_14(.reset(effective_rst), .clk(clk),  .in_a(a9_13to9_14), .in_b(b8_14to9_14),  .out_a(a9_14to9_15), .out_b(b9_14to10_14), .out_c(matrixC9_14));
processing_element pe9_15(.reset(effective_rst), .clk(clk),  .in_a(a9_14to9_15), .in_b(b8_15to9_15),  .out_a(a9_15to9_16), .out_b(b9_15to10_15), .out_c(matrixC9_15));
processing_element pe9_16(.reset(effective_rst), .clk(clk),  .in_a(a9_15to9_16), .in_b(b8_16to9_16),  .out_a(a9_16to9_17), .out_b(b9_16to10_16), .out_c(matrixC9_16));
processing_element pe9_17(.reset(effective_rst), .clk(clk),  .in_a(a9_16to9_17), .in_b(b8_17to9_17),  .out_a(a9_17to9_18), .out_b(b9_17to10_17), .out_c(matrixC9_17));
processing_element pe9_18(.reset(effective_rst), .clk(clk),  .in_a(a9_17to9_18), .in_b(b8_18to9_18),  .out_a(a9_18to9_19), .out_b(b9_18to10_18), .out_c(matrixC9_18));
processing_element pe9_19(.reset(effective_rst), .clk(clk),  .in_a(a9_18to9_19), .in_b(b8_19to9_19),  .out_a(a9_19to9_20), .out_b(b9_19to10_19), .out_c(matrixC9_19));
processing_element pe9_20(.reset(effective_rst), .clk(clk),  .in_a(a9_19to9_20), .in_b(b8_20to9_20),  .out_a(a9_20to9_21), .out_b(b9_20to10_20), .out_c(matrixC9_20));
processing_element pe9_21(.reset(effective_rst), .clk(clk),  .in_a(a9_20to9_21), .in_b(b8_21to9_21),  .out_a(a9_21to9_22), .out_b(b9_21to10_21), .out_c(matrixC9_21));
processing_element pe9_22(.reset(effective_rst), .clk(clk),  .in_a(a9_21to9_22), .in_b(b8_22to9_22),  .out_a(a9_22to9_23), .out_b(b9_22to10_22), .out_c(matrixC9_22));
processing_element pe9_23(.reset(effective_rst), .clk(clk),  .in_a(a9_22to9_23), .in_b(b8_23to9_23),  .out_a(a9_23to9_24), .out_b(b9_23to10_23), .out_c(matrixC9_23));
processing_element pe9_24(.reset(effective_rst), .clk(clk),  .in_a(a9_23to9_24), .in_b(b8_24to9_24),  .out_a(a9_24to9_25), .out_b(b9_24to10_24), .out_c(matrixC9_24));
processing_element pe9_25(.reset(effective_rst), .clk(clk),  .in_a(a9_24to9_25), .in_b(b8_25to9_25),  .out_a(a9_25to9_26), .out_b(b9_25to10_25), .out_c(matrixC9_25));
processing_element pe9_26(.reset(effective_rst), .clk(clk),  .in_a(a9_25to9_26), .in_b(b8_26to9_26),  .out_a(a9_26to9_27), .out_b(b9_26to10_26), .out_c(matrixC9_26));
processing_element pe9_27(.reset(effective_rst), .clk(clk),  .in_a(a9_26to9_27), .in_b(b8_27to9_27),  .out_a(a9_27to9_28), .out_b(b9_27to10_27), .out_c(matrixC9_27));
processing_element pe9_28(.reset(effective_rst), .clk(clk),  .in_a(a9_27to9_28), .in_b(b8_28to9_28),  .out_a(a9_28to9_29), .out_b(b9_28to10_28), .out_c(matrixC9_28));
processing_element pe9_29(.reset(effective_rst), .clk(clk),  .in_a(a9_28to9_29), .in_b(b8_29to9_29),  .out_a(a9_29to9_30), .out_b(b9_29to10_29), .out_c(matrixC9_29));
processing_element pe9_30(.reset(effective_rst), .clk(clk),  .in_a(a9_29to9_30), .in_b(b8_30to9_30),  .out_a(a9_30to9_31), .out_b(b9_30to10_30), .out_c(matrixC9_30));
processing_element pe9_31(.reset(effective_rst), .clk(clk),  .in_a(a9_30to9_31), .in_b(b8_31to9_31),  .out_a(a9_31to9_32), .out_b(b9_31to10_31), .out_c(matrixC9_31));
processing_element pe10_1(.reset(effective_rst), .clk(clk),  .in_a(a10_0to10_1), .in_b(b9_1to10_1),  .out_a(a10_1to10_2), .out_b(b10_1to11_1), .out_c(matrixC10_1));
processing_element pe10_2(.reset(effective_rst), .clk(clk),  .in_a(a10_1to10_2), .in_b(b9_2to10_2),  .out_a(a10_2to10_3), .out_b(b10_2to11_2), .out_c(matrixC10_2));
processing_element pe10_3(.reset(effective_rst), .clk(clk),  .in_a(a10_2to10_3), .in_b(b9_3to10_3),  .out_a(a10_3to10_4), .out_b(b10_3to11_3), .out_c(matrixC10_3));
processing_element pe10_4(.reset(effective_rst), .clk(clk),  .in_a(a10_3to10_4), .in_b(b9_4to10_4),  .out_a(a10_4to10_5), .out_b(b10_4to11_4), .out_c(matrixC10_4));
processing_element pe10_5(.reset(effective_rst), .clk(clk),  .in_a(a10_4to10_5), .in_b(b9_5to10_5),  .out_a(a10_5to10_6), .out_b(b10_5to11_5), .out_c(matrixC10_5));
processing_element pe10_6(.reset(effective_rst), .clk(clk),  .in_a(a10_5to10_6), .in_b(b9_6to10_6),  .out_a(a10_6to10_7), .out_b(b10_6to11_6), .out_c(matrixC10_6));
processing_element pe10_7(.reset(effective_rst), .clk(clk),  .in_a(a10_6to10_7), .in_b(b9_7to10_7),  .out_a(a10_7to10_8), .out_b(b10_7to11_7), .out_c(matrixC10_7));
processing_element pe10_8(.reset(effective_rst), .clk(clk),  .in_a(a10_7to10_8), .in_b(b9_8to10_8),  .out_a(a10_8to10_9), .out_b(b10_8to11_8), .out_c(matrixC10_8));
processing_element pe10_9(.reset(effective_rst), .clk(clk),  .in_a(a10_8to10_9), .in_b(b9_9to10_9),  .out_a(a10_9to10_10), .out_b(b10_9to11_9), .out_c(matrixC10_9));
processing_element pe10_10(.reset(effective_rst), .clk(clk),  .in_a(a10_9to10_10), .in_b(b9_10to10_10),  .out_a(a10_10to10_11), .out_b(b10_10to11_10), .out_c(matrixC10_10));
processing_element pe10_11(.reset(effective_rst), .clk(clk),  .in_a(a10_10to10_11), .in_b(b9_11to10_11),  .out_a(a10_11to10_12), .out_b(b10_11to11_11), .out_c(matrixC10_11));
processing_element pe10_12(.reset(effective_rst), .clk(clk),  .in_a(a10_11to10_12), .in_b(b9_12to10_12),  .out_a(a10_12to10_13), .out_b(b10_12to11_12), .out_c(matrixC10_12));
processing_element pe10_13(.reset(effective_rst), .clk(clk),  .in_a(a10_12to10_13), .in_b(b9_13to10_13),  .out_a(a10_13to10_14), .out_b(b10_13to11_13), .out_c(matrixC10_13));
processing_element pe10_14(.reset(effective_rst), .clk(clk),  .in_a(a10_13to10_14), .in_b(b9_14to10_14),  .out_a(a10_14to10_15), .out_b(b10_14to11_14), .out_c(matrixC10_14));
processing_element pe10_15(.reset(effective_rst), .clk(clk),  .in_a(a10_14to10_15), .in_b(b9_15to10_15),  .out_a(a10_15to10_16), .out_b(b10_15to11_15), .out_c(matrixC10_15));
processing_element pe10_16(.reset(effective_rst), .clk(clk),  .in_a(a10_15to10_16), .in_b(b9_16to10_16),  .out_a(a10_16to10_17), .out_b(b10_16to11_16), .out_c(matrixC10_16));
processing_element pe10_17(.reset(effective_rst), .clk(clk),  .in_a(a10_16to10_17), .in_b(b9_17to10_17),  .out_a(a10_17to10_18), .out_b(b10_17to11_17), .out_c(matrixC10_17));
processing_element pe10_18(.reset(effective_rst), .clk(clk),  .in_a(a10_17to10_18), .in_b(b9_18to10_18),  .out_a(a10_18to10_19), .out_b(b10_18to11_18), .out_c(matrixC10_18));
processing_element pe10_19(.reset(effective_rst), .clk(clk),  .in_a(a10_18to10_19), .in_b(b9_19to10_19),  .out_a(a10_19to10_20), .out_b(b10_19to11_19), .out_c(matrixC10_19));
processing_element pe10_20(.reset(effective_rst), .clk(clk),  .in_a(a10_19to10_20), .in_b(b9_20to10_20),  .out_a(a10_20to10_21), .out_b(b10_20to11_20), .out_c(matrixC10_20));
processing_element pe10_21(.reset(effective_rst), .clk(clk),  .in_a(a10_20to10_21), .in_b(b9_21to10_21),  .out_a(a10_21to10_22), .out_b(b10_21to11_21), .out_c(matrixC10_21));
processing_element pe10_22(.reset(effective_rst), .clk(clk),  .in_a(a10_21to10_22), .in_b(b9_22to10_22),  .out_a(a10_22to10_23), .out_b(b10_22to11_22), .out_c(matrixC10_22));
processing_element pe10_23(.reset(effective_rst), .clk(clk),  .in_a(a10_22to10_23), .in_b(b9_23to10_23),  .out_a(a10_23to10_24), .out_b(b10_23to11_23), .out_c(matrixC10_23));
processing_element pe10_24(.reset(effective_rst), .clk(clk),  .in_a(a10_23to10_24), .in_b(b9_24to10_24),  .out_a(a10_24to10_25), .out_b(b10_24to11_24), .out_c(matrixC10_24));
processing_element pe10_25(.reset(effective_rst), .clk(clk),  .in_a(a10_24to10_25), .in_b(b9_25to10_25),  .out_a(a10_25to10_26), .out_b(b10_25to11_25), .out_c(matrixC10_25));
processing_element pe10_26(.reset(effective_rst), .clk(clk),  .in_a(a10_25to10_26), .in_b(b9_26to10_26),  .out_a(a10_26to10_27), .out_b(b10_26to11_26), .out_c(matrixC10_26));
processing_element pe10_27(.reset(effective_rst), .clk(clk),  .in_a(a10_26to10_27), .in_b(b9_27to10_27),  .out_a(a10_27to10_28), .out_b(b10_27to11_27), .out_c(matrixC10_27));
processing_element pe10_28(.reset(effective_rst), .clk(clk),  .in_a(a10_27to10_28), .in_b(b9_28to10_28),  .out_a(a10_28to10_29), .out_b(b10_28to11_28), .out_c(matrixC10_28));
processing_element pe10_29(.reset(effective_rst), .clk(clk),  .in_a(a10_28to10_29), .in_b(b9_29to10_29),  .out_a(a10_29to10_30), .out_b(b10_29to11_29), .out_c(matrixC10_29));
processing_element pe10_30(.reset(effective_rst), .clk(clk),  .in_a(a10_29to10_30), .in_b(b9_30to10_30),  .out_a(a10_30to10_31), .out_b(b10_30to11_30), .out_c(matrixC10_30));
processing_element pe10_31(.reset(effective_rst), .clk(clk),  .in_a(a10_30to10_31), .in_b(b9_31to10_31),  .out_a(a10_31to10_32), .out_b(b10_31to11_31), .out_c(matrixC10_31));
processing_element pe11_1(.reset(effective_rst), .clk(clk),  .in_a(a11_0to11_1), .in_b(b10_1to11_1),  .out_a(a11_1to11_2), .out_b(b11_1to12_1), .out_c(matrixC11_1));
processing_element pe11_2(.reset(effective_rst), .clk(clk),  .in_a(a11_1to11_2), .in_b(b10_2to11_2),  .out_a(a11_2to11_3), .out_b(b11_2to12_2), .out_c(matrixC11_2));
processing_element pe11_3(.reset(effective_rst), .clk(clk),  .in_a(a11_2to11_3), .in_b(b10_3to11_3),  .out_a(a11_3to11_4), .out_b(b11_3to12_3), .out_c(matrixC11_3));
processing_element pe11_4(.reset(effective_rst), .clk(clk),  .in_a(a11_3to11_4), .in_b(b10_4to11_4),  .out_a(a11_4to11_5), .out_b(b11_4to12_4), .out_c(matrixC11_4));
processing_element pe11_5(.reset(effective_rst), .clk(clk),  .in_a(a11_4to11_5), .in_b(b10_5to11_5),  .out_a(a11_5to11_6), .out_b(b11_5to12_5), .out_c(matrixC11_5));
processing_element pe11_6(.reset(effective_rst), .clk(clk),  .in_a(a11_5to11_6), .in_b(b10_6to11_6),  .out_a(a11_6to11_7), .out_b(b11_6to12_6), .out_c(matrixC11_6));
processing_element pe11_7(.reset(effective_rst), .clk(clk),  .in_a(a11_6to11_7), .in_b(b10_7to11_7),  .out_a(a11_7to11_8), .out_b(b11_7to12_7), .out_c(matrixC11_7));
processing_element pe11_8(.reset(effective_rst), .clk(clk),  .in_a(a11_7to11_8), .in_b(b10_8to11_8),  .out_a(a11_8to11_9), .out_b(b11_8to12_8), .out_c(matrixC11_8));
processing_element pe11_9(.reset(effective_rst), .clk(clk),  .in_a(a11_8to11_9), .in_b(b10_9to11_9),  .out_a(a11_9to11_10), .out_b(b11_9to12_9), .out_c(matrixC11_9));
processing_element pe11_10(.reset(effective_rst), .clk(clk),  .in_a(a11_9to11_10), .in_b(b10_10to11_10),  .out_a(a11_10to11_11), .out_b(b11_10to12_10), .out_c(matrixC11_10));
processing_element pe11_11(.reset(effective_rst), .clk(clk),  .in_a(a11_10to11_11), .in_b(b10_11to11_11),  .out_a(a11_11to11_12), .out_b(b11_11to12_11), .out_c(matrixC11_11));
processing_element pe11_12(.reset(effective_rst), .clk(clk),  .in_a(a11_11to11_12), .in_b(b10_12to11_12),  .out_a(a11_12to11_13), .out_b(b11_12to12_12), .out_c(matrixC11_12));
processing_element pe11_13(.reset(effective_rst), .clk(clk),  .in_a(a11_12to11_13), .in_b(b10_13to11_13),  .out_a(a11_13to11_14), .out_b(b11_13to12_13), .out_c(matrixC11_13));
processing_element pe11_14(.reset(effective_rst), .clk(clk),  .in_a(a11_13to11_14), .in_b(b10_14to11_14),  .out_a(a11_14to11_15), .out_b(b11_14to12_14), .out_c(matrixC11_14));
processing_element pe11_15(.reset(effective_rst), .clk(clk),  .in_a(a11_14to11_15), .in_b(b10_15to11_15),  .out_a(a11_15to11_16), .out_b(b11_15to12_15), .out_c(matrixC11_15));
processing_element pe11_16(.reset(effective_rst), .clk(clk),  .in_a(a11_15to11_16), .in_b(b10_16to11_16),  .out_a(a11_16to11_17), .out_b(b11_16to12_16), .out_c(matrixC11_16));
processing_element pe11_17(.reset(effective_rst), .clk(clk),  .in_a(a11_16to11_17), .in_b(b10_17to11_17),  .out_a(a11_17to11_18), .out_b(b11_17to12_17), .out_c(matrixC11_17));
processing_element pe11_18(.reset(effective_rst), .clk(clk),  .in_a(a11_17to11_18), .in_b(b10_18to11_18),  .out_a(a11_18to11_19), .out_b(b11_18to12_18), .out_c(matrixC11_18));
processing_element pe11_19(.reset(effective_rst), .clk(clk),  .in_a(a11_18to11_19), .in_b(b10_19to11_19),  .out_a(a11_19to11_20), .out_b(b11_19to12_19), .out_c(matrixC11_19));
processing_element pe11_20(.reset(effective_rst), .clk(clk),  .in_a(a11_19to11_20), .in_b(b10_20to11_20),  .out_a(a11_20to11_21), .out_b(b11_20to12_20), .out_c(matrixC11_20));
processing_element pe11_21(.reset(effective_rst), .clk(clk),  .in_a(a11_20to11_21), .in_b(b10_21to11_21),  .out_a(a11_21to11_22), .out_b(b11_21to12_21), .out_c(matrixC11_21));
processing_element pe11_22(.reset(effective_rst), .clk(clk),  .in_a(a11_21to11_22), .in_b(b10_22to11_22),  .out_a(a11_22to11_23), .out_b(b11_22to12_22), .out_c(matrixC11_22));
processing_element pe11_23(.reset(effective_rst), .clk(clk),  .in_a(a11_22to11_23), .in_b(b10_23to11_23),  .out_a(a11_23to11_24), .out_b(b11_23to12_23), .out_c(matrixC11_23));
processing_element pe11_24(.reset(effective_rst), .clk(clk),  .in_a(a11_23to11_24), .in_b(b10_24to11_24),  .out_a(a11_24to11_25), .out_b(b11_24to12_24), .out_c(matrixC11_24));
processing_element pe11_25(.reset(effective_rst), .clk(clk),  .in_a(a11_24to11_25), .in_b(b10_25to11_25),  .out_a(a11_25to11_26), .out_b(b11_25to12_25), .out_c(matrixC11_25));
processing_element pe11_26(.reset(effective_rst), .clk(clk),  .in_a(a11_25to11_26), .in_b(b10_26to11_26),  .out_a(a11_26to11_27), .out_b(b11_26to12_26), .out_c(matrixC11_26));
processing_element pe11_27(.reset(effective_rst), .clk(clk),  .in_a(a11_26to11_27), .in_b(b10_27to11_27),  .out_a(a11_27to11_28), .out_b(b11_27to12_27), .out_c(matrixC11_27));
processing_element pe11_28(.reset(effective_rst), .clk(clk),  .in_a(a11_27to11_28), .in_b(b10_28to11_28),  .out_a(a11_28to11_29), .out_b(b11_28to12_28), .out_c(matrixC11_28));
processing_element pe11_29(.reset(effective_rst), .clk(clk),  .in_a(a11_28to11_29), .in_b(b10_29to11_29),  .out_a(a11_29to11_30), .out_b(b11_29to12_29), .out_c(matrixC11_29));
processing_element pe11_30(.reset(effective_rst), .clk(clk),  .in_a(a11_29to11_30), .in_b(b10_30to11_30),  .out_a(a11_30to11_31), .out_b(b11_30to12_30), .out_c(matrixC11_30));
processing_element pe11_31(.reset(effective_rst), .clk(clk),  .in_a(a11_30to11_31), .in_b(b10_31to11_31),  .out_a(a11_31to11_32), .out_b(b11_31to12_31), .out_c(matrixC11_31));
processing_element pe12_1(.reset(effective_rst), .clk(clk),  .in_a(a12_0to12_1), .in_b(b11_1to12_1),  .out_a(a12_1to12_2), .out_b(b12_1to13_1), .out_c(matrixC12_1));
processing_element pe12_2(.reset(effective_rst), .clk(clk),  .in_a(a12_1to12_2), .in_b(b11_2to12_2),  .out_a(a12_2to12_3), .out_b(b12_2to13_2), .out_c(matrixC12_2));
processing_element pe12_3(.reset(effective_rst), .clk(clk),  .in_a(a12_2to12_3), .in_b(b11_3to12_3),  .out_a(a12_3to12_4), .out_b(b12_3to13_3), .out_c(matrixC12_3));
processing_element pe12_4(.reset(effective_rst), .clk(clk),  .in_a(a12_3to12_4), .in_b(b11_4to12_4),  .out_a(a12_4to12_5), .out_b(b12_4to13_4), .out_c(matrixC12_4));
processing_element pe12_5(.reset(effective_rst), .clk(clk),  .in_a(a12_4to12_5), .in_b(b11_5to12_5),  .out_a(a12_5to12_6), .out_b(b12_5to13_5), .out_c(matrixC12_5));
processing_element pe12_6(.reset(effective_rst), .clk(clk),  .in_a(a12_5to12_6), .in_b(b11_6to12_6),  .out_a(a12_6to12_7), .out_b(b12_6to13_6), .out_c(matrixC12_6));
processing_element pe12_7(.reset(effective_rst), .clk(clk),  .in_a(a12_6to12_7), .in_b(b11_7to12_7),  .out_a(a12_7to12_8), .out_b(b12_7to13_7), .out_c(matrixC12_7));
processing_element pe12_8(.reset(effective_rst), .clk(clk),  .in_a(a12_7to12_8), .in_b(b11_8to12_8),  .out_a(a12_8to12_9), .out_b(b12_8to13_8), .out_c(matrixC12_8));
processing_element pe12_9(.reset(effective_rst), .clk(clk),  .in_a(a12_8to12_9), .in_b(b11_9to12_9),  .out_a(a12_9to12_10), .out_b(b12_9to13_9), .out_c(matrixC12_9));
processing_element pe12_10(.reset(effective_rst), .clk(clk),  .in_a(a12_9to12_10), .in_b(b11_10to12_10),  .out_a(a12_10to12_11), .out_b(b12_10to13_10), .out_c(matrixC12_10));
processing_element pe12_11(.reset(effective_rst), .clk(clk),  .in_a(a12_10to12_11), .in_b(b11_11to12_11),  .out_a(a12_11to12_12), .out_b(b12_11to13_11), .out_c(matrixC12_11));
processing_element pe12_12(.reset(effective_rst), .clk(clk),  .in_a(a12_11to12_12), .in_b(b11_12to12_12),  .out_a(a12_12to12_13), .out_b(b12_12to13_12), .out_c(matrixC12_12));
processing_element pe12_13(.reset(effective_rst), .clk(clk),  .in_a(a12_12to12_13), .in_b(b11_13to12_13),  .out_a(a12_13to12_14), .out_b(b12_13to13_13), .out_c(matrixC12_13));
processing_element pe12_14(.reset(effective_rst), .clk(clk),  .in_a(a12_13to12_14), .in_b(b11_14to12_14),  .out_a(a12_14to12_15), .out_b(b12_14to13_14), .out_c(matrixC12_14));
processing_element pe12_15(.reset(effective_rst), .clk(clk),  .in_a(a12_14to12_15), .in_b(b11_15to12_15),  .out_a(a12_15to12_16), .out_b(b12_15to13_15), .out_c(matrixC12_15));
processing_element pe12_16(.reset(effective_rst), .clk(clk),  .in_a(a12_15to12_16), .in_b(b11_16to12_16),  .out_a(a12_16to12_17), .out_b(b12_16to13_16), .out_c(matrixC12_16));
processing_element pe12_17(.reset(effective_rst), .clk(clk),  .in_a(a12_16to12_17), .in_b(b11_17to12_17),  .out_a(a12_17to12_18), .out_b(b12_17to13_17), .out_c(matrixC12_17));
processing_element pe12_18(.reset(effective_rst), .clk(clk),  .in_a(a12_17to12_18), .in_b(b11_18to12_18),  .out_a(a12_18to12_19), .out_b(b12_18to13_18), .out_c(matrixC12_18));
processing_element pe12_19(.reset(effective_rst), .clk(clk),  .in_a(a12_18to12_19), .in_b(b11_19to12_19),  .out_a(a12_19to12_20), .out_b(b12_19to13_19), .out_c(matrixC12_19));
processing_element pe12_20(.reset(effective_rst), .clk(clk),  .in_a(a12_19to12_20), .in_b(b11_20to12_20),  .out_a(a12_20to12_21), .out_b(b12_20to13_20), .out_c(matrixC12_20));
processing_element pe12_21(.reset(effective_rst), .clk(clk),  .in_a(a12_20to12_21), .in_b(b11_21to12_21),  .out_a(a12_21to12_22), .out_b(b12_21to13_21), .out_c(matrixC12_21));
processing_element pe12_22(.reset(effective_rst), .clk(clk),  .in_a(a12_21to12_22), .in_b(b11_22to12_22),  .out_a(a12_22to12_23), .out_b(b12_22to13_22), .out_c(matrixC12_22));
processing_element pe12_23(.reset(effective_rst), .clk(clk),  .in_a(a12_22to12_23), .in_b(b11_23to12_23),  .out_a(a12_23to12_24), .out_b(b12_23to13_23), .out_c(matrixC12_23));
processing_element pe12_24(.reset(effective_rst), .clk(clk),  .in_a(a12_23to12_24), .in_b(b11_24to12_24),  .out_a(a12_24to12_25), .out_b(b12_24to13_24), .out_c(matrixC12_24));
processing_element pe12_25(.reset(effective_rst), .clk(clk),  .in_a(a12_24to12_25), .in_b(b11_25to12_25),  .out_a(a12_25to12_26), .out_b(b12_25to13_25), .out_c(matrixC12_25));
processing_element pe12_26(.reset(effective_rst), .clk(clk),  .in_a(a12_25to12_26), .in_b(b11_26to12_26),  .out_a(a12_26to12_27), .out_b(b12_26to13_26), .out_c(matrixC12_26));
processing_element pe12_27(.reset(effective_rst), .clk(clk),  .in_a(a12_26to12_27), .in_b(b11_27to12_27),  .out_a(a12_27to12_28), .out_b(b12_27to13_27), .out_c(matrixC12_27));
processing_element pe12_28(.reset(effective_rst), .clk(clk),  .in_a(a12_27to12_28), .in_b(b11_28to12_28),  .out_a(a12_28to12_29), .out_b(b12_28to13_28), .out_c(matrixC12_28));
processing_element pe12_29(.reset(effective_rst), .clk(clk),  .in_a(a12_28to12_29), .in_b(b11_29to12_29),  .out_a(a12_29to12_30), .out_b(b12_29to13_29), .out_c(matrixC12_29));
processing_element pe12_30(.reset(effective_rst), .clk(clk),  .in_a(a12_29to12_30), .in_b(b11_30to12_30),  .out_a(a12_30to12_31), .out_b(b12_30to13_30), .out_c(matrixC12_30));
processing_element pe12_31(.reset(effective_rst), .clk(clk),  .in_a(a12_30to12_31), .in_b(b11_31to12_31),  .out_a(a12_31to12_32), .out_b(b12_31to13_31), .out_c(matrixC12_31));
processing_element pe13_1(.reset(effective_rst), .clk(clk),  .in_a(a13_0to13_1), .in_b(b12_1to13_1),  .out_a(a13_1to13_2), .out_b(b13_1to14_1), .out_c(matrixC13_1));
processing_element pe13_2(.reset(effective_rst), .clk(clk),  .in_a(a13_1to13_2), .in_b(b12_2to13_2),  .out_a(a13_2to13_3), .out_b(b13_2to14_2), .out_c(matrixC13_2));
processing_element pe13_3(.reset(effective_rst), .clk(clk),  .in_a(a13_2to13_3), .in_b(b12_3to13_3),  .out_a(a13_3to13_4), .out_b(b13_3to14_3), .out_c(matrixC13_3));
processing_element pe13_4(.reset(effective_rst), .clk(clk),  .in_a(a13_3to13_4), .in_b(b12_4to13_4),  .out_a(a13_4to13_5), .out_b(b13_4to14_4), .out_c(matrixC13_4));
processing_element pe13_5(.reset(effective_rst), .clk(clk),  .in_a(a13_4to13_5), .in_b(b12_5to13_5),  .out_a(a13_5to13_6), .out_b(b13_5to14_5), .out_c(matrixC13_5));
processing_element pe13_6(.reset(effective_rst), .clk(clk),  .in_a(a13_5to13_6), .in_b(b12_6to13_6),  .out_a(a13_6to13_7), .out_b(b13_6to14_6), .out_c(matrixC13_6));
processing_element pe13_7(.reset(effective_rst), .clk(clk),  .in_a(a13_6to13_7), .in_b(b12_7to13_7),  .out_a(a13_7to13_8), .out_b(b13_7to14_7), .out_c(matrixC13_7));
processing_element pe13_8(.reset(effective_rst), .clk(clk),  .in_a(a13_7to13_8), .in_b(b12_8to13_8),  .out_a(a13_8to13_9), .out_b(b13_8to14_8), .out_c(matrixC13_8));
processing_element pe13_9(.reset(effective_rst), .clk(clk),  .in_a(a13_8to13_9), .in_b(b12_9to13_9),  .out_a(a13_9to13_10), .out_b(b13_9to14_9), .out_c(matrixC13_9));
processing_element pe13_10(.reset(effective_rst), .clk(clk),  .in_a(a13_9to13_10), .in_b(b12_10to13_10),  .out_a(a13_10to13_11), .out_b(b13_10to14_10), .out_c(matrixC13_10));
processing_element pe13_11(.reset(effective_rst), .clk(clk),  .in_a(a13_10to13_11), .in_b(b12_11to13_11),  .out_a(a13_11to13_12), .out_b(b13_11to14_11), .out_c(matrixC13_11));
processing_element pe13_12(.reset(effective_rst), .clk(clk),  .in_a(a13_11to13_12), .in_b(b12_12to13_12),  .out_a(a13_12to13_13), .out_b(b13_12to14_12), .out_c(matrixC13_12));
processing_element pe13_13(.reset(effective_rst), .clk(clk),  .in_a(a13_12to13_13), .in_b(b12_13to13_13),  .out_a(a13_13to13_14), .out_b(b13_13to14_13), .out_c(matrixC13_13));
processing_element pe13_14(.reset(effective_rst), .clk(clk),  .in_a(a13_13to13_14), .in_b(b12_14to13_14),  .out_a(a13_14to13_15), .out_b(b13_14to14_14), .out_c(matrixC13_14));
processing_element pe13_15(.reset(effective_rst), .clk(clk),  .in_a(a13_14to13_15), .in_b(b12_15to13_15),  .out_a(a13_15to13_16), .out_b(b13_15to14_15), .out_c(matrixC13_15));
processing_element pe13_16(.reset(effective_rst), .clk(clk),  .in_a(a13_15to13_16), .in_b(b12_16to13_16),  .out_a(a13_16to13_17), .out_b(b13_16to14_16), .out_c(matrixC13_16));
processing_element pe13_17(.reset(effective_rst), .clk(clk),  .in_a(a13_16to13_17), .in_b(b12_17to13_17),  .out_a(a13_17to13_18), .out_b(b13_17to14_17), .out_c(matrixC13_17));
processing_element pe13_18(.reset(effective_rst), .clk(clk),  .in_a(a13_17to13_18), .in_b(b12_18to13_18),  .out_a(a13_18to13_19), .out_b(b13_18to14_18), .out_c(matrixC13_18));
processing_element pe13_19(.reset(effective_rst), .clk(clk),  .in_a(a13_18to13_19), .in_b(b12_19to13_19),  .out_a(a13_19to13_20), .out_b(b13_19to14_19), .out_c(matrixC13_19));
processing_element pe13_20(.reset(effective_rst), .clk(clk),  .in_a(a13_19to13_20), .in_b(b12_20to13_20),  .out_a(a13_20to13_21), .out_b(b13_20to14_20), .out_c(matrixC13_20));
processing_element pe13_21(.reset(effective_rst), .clk(clk),  .in_a(a13_20to13_21), .in_b(b12_21to13_21),  .out_a(a13_21to13_22), .out_b(b13_21to14_21), .out_c(matrixC13_21));
processing_element pe13_22(.reset(effective_rst), .clk(clk),  .in_a(a13_21to13_22), .in_b(b12_22to13_22),  .out_a(a13_22to13_23), .out_b(b13_22to14_22), .out_c(matrixC13_22));
processing_element pe13_23(.reset(effective_rst), .clk(clk),  .in_a(a13_22to13_23), .in_b(b12_23to13_23),  .out_a(a13_23to13_24), .out_b(b13_23to14_23), .out_c(matrixC13_23));
processing_element pe13_24(.reset(effective_rst), .clk(clk),  .in_a(a13_23to13_24), .in_b(b12_24to13_24),  .out_a(a13_24to13_25), .out_b(b13_24to14_24), .out_c(matrixC13_24));
processing_element pe13_25(.reset(effective_rst), .clk(clk),  .in_a(a13_24to13_25), .in_b(b12_25to13_25),  .out_a(a13_25to13_26), .out_b(b13_25to14_25), .out_c(matrixC13_25));
processing_element pe13_26(.reset(effective_rst), .clk(clk),  .in_a(a13_25to13_26), .in_b(b12_26to13_26),  .out_a(a13_26to13_27), .out_b(b13_26to14_26), .out_c(matrixC13_26));
processing_element pe13_27(.reset(effective_rst), .clk(clk),  .in_a(a13_26to13_27), .in_b(b12_27to13_27),  .out_a(a13_27to13_28), .out_b(b13_27to14_27), .out_c(matrixC13_27));
processing_element pe13_28(.reset(effective_rst), .clk(clk),  .in_a(a13_27to13_28), .in_b(b12_28to13_28),  .out_a(a13_28to13_29), .out_b(b13_28to14_28), .out_c(matrixC13_28));
processing_element pe13_29(.reset(effective_rst), .clk(clk),  .in_a(a13_28to13_29), .in_b(b12_29to13_29),  .out_a(a13_29to13_30), .out_b(b13_29to14_29), .out_c(matrixC13_29));
processing_element pe13_30(.reset(effective_rst), .clk(clk),  .in_a(a13_29to13_30), .in_b(b12_30to13_30),  .out_a(a13_30to13_31), .out_b(b13_30to14_30), .out_c(matrixC13_30));
processing_element pe13_31(.reset(effective_rst), .clk(clk),  .in_a(a13_30to13_31), .in_b(b12_31to13_31),  .out_a(a13_31to13_32), .out_b(b13_31to14_31), .out_c(matrixC13_31));
processing_element pe14_1(.reset(effective_rst), .clk(clk),  .in_a(a14_0to14_1), .in_b(b13_1to14_1),  .out_a(a14_1to14_2), .out_b(b14_1to15_1), .out_c(matrixC14_1));
processing_element pe14_2(.reset(effective_rst), .clk(clk),  .in_a(a14_1to14_2), .in_b(b13_2to14_2),  .out_a(a14_2to14_3), .out_b(b14_2to15_2), .out_c(matrixC14_2));
processing_element pe14_3(.reset(effective_rst), .clk(clk),  .in_a(a14_2to14_3), .in_b(b13_3to14_3),  .out_a(a14_3to14_4), .out_b(b14_3to15_3), .out_c(matrixC14_3));
processing_element pe14_4(.reset(effective_rst), .clk(clk),  .in_a(a14_3to14_4), .in_b(b13_4to14_4),  .out_a(a14_4to14_5), .out_b(b14_4to15_4), .out_c(matrixC14_4));
processing_element pe14_5(.reset(effective_rst), .clk(clk),  .in_a(a14_4to14_5), .in_b(b13_5to14_5),  .out_a(a14_5to14_6), .out_b(b14_5to15_5), .out_c(matrixC14_5));
processing_element pe14_6(.reset(effective_rst), .clk(clk),  .in_a(a14_5to14_6), .in_b(b13_6to14_6),  .out_a(a14_6to14_7), .out_b(b14_6to15_6), .out_c(matrixC14_6));
processing_element pe14_7(.reset(effective_rst), .clk(clk),  .in_a(a14_6to14_7), .in_b(b13_7to14_7),  .out_a(a14_7to14_8), .out_b(b14_7to15_7), .out_c(matrixC14_7));
processing_element pe14_8(.reset(effective_rst), .clk(clk),  .in_a(a14_7to14_8), .in_b(b13_8to14_8),  .out_a(a14_8to14_9), .out_b(b14_8to15_8), .out_c(matrixC14_8));
processing_element pe14_9(.reset(effective_rst), .clk(clk),  .in_a(a14_8to14_9), .in_b(b13_9to14_9),  .out_a(a14_9to14_10), .out_b(b14_9to15_9), .out_c(matrixC14_9));
processing_element pe14_10(.reset(effective_rst), .clk(clk),  .in_a(a14_9to14_10), .in_b(b13_10to14_10),  .out_a(a14_10to14_11), .out_b(b14_10to15_10), .out_c(matrixC14_10));
processing_element pe14_11(.reset(effective_rst), .clk(clk),  .in_a(a14_10to14_11), .in_b(b13_11to14_11),  .out_a(a14_11to14_12), .out_b(b14_11to15_11), .out_c(matrixC14_11));
processing_element pe14_12(.reset(effective_rst), .clk(clk),  .in_a(a14_11to14_12), .in_b(b13_12to14_12),  .out_a(a14_12to14_13), .out_b(b14_12to15_12), .out_c(matrixC14_12));
processing_element pe14_13(.reset(effective_rst), .clk(clk),  .in_a(a14_12to14_13), .in_b(b13_13to14_13),  .out_a(a14_13to14_14), .out_b(b14_13to15_13), .out_c(matrixC14_13));
processing_element pe14_14(.reset(effective_rst), .clk(clk),  .in_a(a14_13to14_14), .in_b(b13_14to14_14),  .out_a(a14_14to14_15), .out_b(b14_14to15_14), .out_c(matrixC14_14));
processing_element pe14_15(.reset(effective_rst), .clk(clk),  .in_a(a14_14to14_15), .in_b(b13_15to14_15),  .out_a(a14_15to14_16), .out_b(b14_15to15_15), .out_c(matrixC14_15));
processing_element pe14_16(.reset(effective_rst), .clk(clk),  .in_a(a14_15to14_16), .in_b(b13_16to14_16),  .out_a(a14_16to14_17), .out_b(b14_16to15_16), .out_c(matrixC14_16));
processing_element pe14_17(.reset(effective_rst), .clk(clk),  .in_a(a14_16to14_17), .in_b(b13_17to14_17),  .out_a(a14_17to14_18), .out_b(b14_17to15_17), .out_c(matrixC14_17));
processing_element pe14_18(.reset(effective_rst), .clk(clk),  .in_a(a14_17to14_18), .in_b(b13_18to14_18),  .out_a(a14_18to14_19), .out_b(b14_18to15_18), .out_c(matrixC14_18));
processing_element pe14_19(.reset(effective_rst), .clk(clk),  .in_a(a14_18to14_19), .in_b(b13_19to14_19),  .out_a(a14_19to14_20), .out_b(b14_19to15_19), .out_c(matrixC14_19));
processing_element pe14_20(.reset(effective_rst), .clk(clk),  .in_a(a14_19to14_20), .in_b(b13_20to14_20),  .out_a(a14_20to14_21), .out_b(b14_20to15_20), .out_c(matrixC14_20));
processing_element pe14_21(.reset(effective_rst), .clk(clk),  .in_a(a14_20to14_21), .in_b(b13_21to14_21),  .out_a(a14_21to14_22), .out_b(b14_21to15_21), .out_c(matrixC14_21));
processing_element pe14_22(.reset(effective_rst), .clk(clk),  .in_a(a14_21to14_22), .in_b(b13_22to14_22),  .out_a(a14_22to14_23), .out_b(b14_22to15_22), .out_c(matrixC14_22));
processing_element pe14_23(.reset(effective_rst), .clk(clk),  .in_a(a14_22to14_23), .in_b(b13_23to14_23),  .out_a(a14_23to14_24), .out_b(b14_23to15_23), .out_c(matrixC14_23));
processing_element pe14_24(.reset(effective_rst), .clk(clk),  .in_a(a14_23to14_24), .in_b(b13_24to14_24),  .out_a(a14_24to14_25), .out_b(b14_24to15_24), .out_c(matrixC14_24));
processing_element pe14_25(.reset(effective_rst), .clk(clk),  .in_a(a14_24to14_25), .in_b(b13_25to14_25),  .out_a(a14_25to14_26), .out_b(b14_25to15_25), .out_c(matrixC14_25));
processing_element pe14_26(.reset(effective_rst), .clk(clk),  .in_a(a14_25to14_26), .in_b(b13_26to14_26),  .out_a(a14_26to14_27), .out_b(b14_26to15_26), .out_c(matrixC14_26));
processing_element pe14_27(.reset(effective_rst), .clk(clk),  .in_a(a14_26to14_27), .in_b(b13_27to14_27),  .out_a(a14_27to14_28), .out_b(b14_27to15_27), .out_c(matrixC14_27));
processing_element pe14_28(.reset(effective_rst), .clk(clk),  .in_a(a14_27to14_28), .in_b(b13_28to14_28),  .out_a(a14_28to14_29), .out_b(b14_28to15_28), .out_c(matrixC14_28));
processing_element pe14_29(.reset(effective_rst), .clk(clk),  .in_a(a14_28to14_29), .in_b(b13_29to14_29),  .out_a(a14_29to14_30), .out_b(b14_29to15_29), .out_c(matrixC14_29));
processing_element pe14_30(.reset(effective_rst), .clk(clk),  .in_a(a14_29to14_30), .in_b(b13_30to14_30),  .out_a(a14_30to14_31), .out_b(b14_30to15_30), .out_c(matrixC14_30));
processing_element pe14_31(.reset(effective_rst), .clk(clk),  .in_a(a14_30to14_31), .in_b(b13_31to14_31),  .out_a(a14_31to14_32), .out_b(b14_31to15_31), .out_c(matrixC14_31));
processing_element pe15_1(.reset(effective_rst), .clk(clk),  .in_a(a15_0to15_1), .in_b(b14_1to15_1),  .out_a(a15_1to15_2), .out_b(b15_1to16_1), .out_c(matrixC15_1));
processing_element pe15_2(.reset(effective_rst), .clk(clk),  .in_a(a15_1to15_2), .in_b(b14_2to15_2),  .out_a(a15_2to15_3), .out_b(b15_2to16_2), .out_c(matrixC15_2));
processing_element pe15_3(.reset(effective_rst), .clk(clk),  .in_a(a15_2to15_3), .in_b(b14_3to15_3),  .out_a(a15_3to15_4), .out_b(b15_3to16_3), .out_c(matrixC15_3));
processing_element pe15_4(.reset(effective_rst), .clk(clk),  .in_a(a15_3to15_4), .in_b(b14_4to15_4),  .out_a(a15_4to15_5), .out_b(b15_4to16_4), .out_c(matrixC15_4));
processing_element pe15_5(.reset(effective_rst), .clk(clk),  .in_a(a15_4to15_5), .in_b(b14_5to15_5),  .out_a(a15_5to15_6), .out_b(b15_5to16_5), .out_c(matrixC15_5));
processing_element pe15_6(.reset(effective_rst), .clk(clk),  .in_a(a15_5to15_6), .in_b(b14_6to15_6),  .out_a(a15_6to15_7), .out_b(b15_6to16_6), .out_c(matrixC15_6));
processing_element pe15_7(.reset(effective_rst), .clk(clk),  .in_a(a15_6to15_7), .in_b(b14_7to15_7),  .out_a(a15_7to15_8), .out_b(b15_7to16_7), .out_c(matrixC15_7));
processing_element pe15_8(.reset(effective_rst), .clk(clk),  .in_a(a15_7to15_8), .in_b(b14_8to15_8),  .out_a(a15_8to15_9), .out_b(b15_8to16_8), .out_c(matrixC15_8));
processing_element pe15_9(.reset(effective_rst), .clk(clk),  .in_a(a15_8to15_9), .in_b(b14_9to15_9),  .out_a(a15_9to15_10), .out_b(b15_9to16_9), .out_c(matrixC15_9));
processing_element pe15_10(.reset(effective_rst), .clk(clk),  .in_a(a15_9to15_10), .in_b(b14_10to15_10),  .out_a(a15_10to15_11), .out_b(b15_10to16_10), .out_c(matrixC15_10));
processing_element pe15_11(.reset(effective_rst), .clk(clk),  .in_a(a15_10to15_11), .in_b(b14_11to15_11),  .out_a(a15_11to15_12), .out_b(b15_11to16_11), .out_c(matrixC15_11));
processing_element pe15_12(.reset(effective_rst), .clk(clk),  .in_a(a15_11to15_12), .in_b(b14_12to15_12),  .out_a(a15_12to15_13), .out_b(b15_12to16_12), .out_c(matrixC15_12));
processing_element pe15_13(.reset(effective_rst), .clk(clk),  .in_a(a15_12to15_13), .in_b(b14_13to15_13),  .out_a(a15_13to15_14), .out_b(b15_13to16_13), .out_c(matrixC15_13));
processing_element pe15_14(.reset(effective_rst), .clk(clk),  .in_a(a15_13to15_14), .in_b(b14_14to15_14),  .out_a(a15_14to15_15), .out_b(b15_14to16_14), .out_c(matrixC15_14));
processing_element pe15_15(.reset(effective_rst), .clk(clk),  .in_a(a15_14to15_15), .in_b(b14_15to15_15),  .out_a(a15_15to15_16), .out_b(b15_15to16_15), .out_c(matrixC15_15));
processing_element pe15_16(.reset(effective_rst), .clk(clk),  .in_a(a15_15to15_16), .in_b(b14_16to15_16),  .out_a(a15_16to15_17), .out_b(b15_16to16_16), .out_c(matrixC15_16));
processing_element pe15_17(.reset(effective_rst), .clk(clk),  .in_a(a15_16to15_17), .in_b(b14_17to15_17),  .out_a(a15_17to15_18), .out_b(b15_17to16_17), .out_c(matrixC15_17));
processing_element pe15_18(.reset(effective_rst), .clk(clk),  .in_a(a15_17to15_18), .in_b(b14_18to15_18),  .out_a(a15_18to15_19), .out_b(b15_18to16_18), .out_c(matrixC15_18));
processing_element pe15_19(.reset(effective_rst), .clk(clk),  .in_a(a15_18to15_19), .in_b(b14_19to15_19),  .out_a(a15_19to15_20), .out_b(b15_19to16_19), .out_c(matrixC15_19));
processing_element pe15_20(.reset(effective_rst), .clk(clk),  .in_a(a15_19to15_20), .in_b(b14_20to15_20),  .out_a(a15_20to15_21), .out_b(b15_20to16_20), .out_c(matrixC15_20));
processing_element pe15_21(.reset(effective_rst), .clk(clk),  .in_a(a15_20to15_21), .in_b(b14_21to15_21),  .out_a(a15_21to15_22), .out_b(b15_21to16_21), .out_c(matrixC15_21));
processing_element pe15_22(.reset(effective_rst), .clk(clk),  .in_a(a15_21to15_22), .in_b(b14_22to15_22),  .out_a(a15_22to15_23), .out_b(b15_22to16_22), .out_c(matrixC15_22));
processing_element pe15_23(.reset(effective_rst), .clk(clk),  .in_a(a15_22to15_23), .in_b(b14_23to15_23),  .out_a(a15_23to15_24), .out_b(b15_23to16_23), .out_c(matrixC15_23));
processing_element pe15_24(.reset(effective_rst), .clk(clk),  .in_a(a15_23to15_24), .in_b(b14_24to15_24),  .out_a(a15_24to15_25), .out_b(b15_24to16_24), .out_c(matrixC15_24));
processing_element pe15_25(.reset(effective_rst), .clk(clk),  .in_a(a15_24to15_25), .in_b(b14_25to15_25),  .out_a(a15_25to15_26), .out_b(b15_25to16_25), .out_c(matrixC15_25));
processing_element pe15_26(.reset(effective_rst), .clk(clk),  .in_a(a15_25to15_26), .in_b(b14_26to15_26),  .out_a(a15_26to15_27), .out_b(b15_26to16_26), .out_c(matrixC15_26));
processing_element pe15_27(.reset(effective_rst), .clk(clk),  .in_a(a15_26to15_27), .in_b(b14_27to15_27),  .out_a(a15_27to15_28), .out_b(b15_27to16_27), .out_c(matrixC15_27));
processing_element pe15_28(.reset(effective_rst), .clk(clk),  .in_a(a15_27to15_28), .in_b(b14_28to15_28),  .out_a(a15_28to15_29), .out_b(b15_28to16_28), .out_c(matrixC15_28));
processing_element pe15_29(.reset(effective_rst), .clk(clk),  .in_a(a15_28to15_29), .in_b(b14_29to15_29),  .out_a(a15_29to15_30), .out_b(b15_29to16_29), .out_c(matrixC15_29));
processing_element pe15_30(.reset(effective_rst), .clk(clk),  .in_a(a15_29to15_30), .in_b(b14_30to15_30),  .out_a(a15_30to15_31), .out_b(b15_30to16_30), .out_c(matrixC15_30));
processing_element pe15_31(.reset(effective_rst), .clk(clk),  .in_a(a15_30to15_31), .in_b(b14_31to15_31),  .out_a(a15_31to15_32), .out_b(b15_31to16_31), .out_c(matrixC15_31));
processing_element pe16_1(.reset(effective_rst), .clk(clk),  .in_a(a16_0to16_1), .in_b(b15_1to16_1),  .out_a(a16_1to16_2), .out_b(b16_1to17_1), .out_c(matrixC16_1));
processing_element pe16_2(.reset(effective_rst), .clk(clk),  .in_a(a16_1to16_2), .in_b(b15_2to16_2),  .out_a(a16_2to16_3), .out_b(b16_2to17_2), .out_c(matrixC16_2));
processing_element pe16_3(.reset(effective_rst), .clk(clk),  .in_a(a16_2to16_3), .in_b(b15_3to16_3),  .out_a(a16_3to16_4), .out_b(b16_3to17_3), .out_c(matrixC16_3));
processing_element pe16_4(.reset(effective_rst), .clk(clk),  .in_a(a16_3to16_4), .in_b(b15_4to16_4),  .out_a(a16_4to16_5), .out_b(b16_4to17_4), .out_c(matrixC16_4));
processing_element pe16_5(.reset(effective_rst), .clk(clk),  .in_a(a16_4to16_5), .in_b(b15_5to16_5),  .out_a(a16_5to16_6), .out_b(b16_5to17_5), .out_c(matrixC16_5));
processing_element pe16_6(.reset(effective_rst), .clk(clk),  .in_a(a16_5to16_6), .in_b(b15_6to16_6),  .out_a(a16_6to16_7), .out_b(b16_6to17_6), .out_c(matrixC16_6));
processing_element pe16_7(.reset(effective_rst), .clk(clk),  .in_a(a16_6to16_7), .in_b(b15_7to16_7),  .out_a(a16_7to16_8), .out_b(b16_7to17_7), .out_c(matrixC16_7));
processing_element pe16_8(.reset(effective_rst), .clk(clk),  .in_a(a16_7to16_8), .in_b(b15_8to16_8),  .out_a(a16_8to16_9), .out_b(b16_8to17_8), .out_c(matrixC16_8));
processing_element pe16_9(.reset(effective_rst), .clk(clk),  .in_a(a16_8to16_9), .in_b(b15_9to16_9),  .out_a(a16_9to16_10), .out_b(b16_9to17_9), .out_c(matrixC16_9));
processing_element pe16_10(.reset(effective_rst), .clk(clk),  .in_a(a16_9to16_10), .in_b(b15_10to16_10),  .out_a(a16_10to16_11), .out_b(b16_10to17_10), .out_c(matrixC16_10));
processing_element pe16_11(.reset(effective_rst), .clk(clk),  .in_a(a16_10to16_11), .in_b(b15_11to16_11),  .out_a(a16_11to16_12), .out_b(b16_11to17_11), .out_c(matrixC16_11));
processing_element pe16_12(.reset(effective_rst), .clk(clk),  .in_a(a16_11to16_12), .in_b(b15_12to16_12),  .out_a(a16_12to16_13), .out_b(b16_12to17_12), .out_c(matrixC16_12));
processing_element pe16_13(.reset(effective_rst), .clk(clk),  .in_a(a16_12to16_13), .in_b(b15_13to16_13),  .out_a(a16_13to16_14), .out_b(b16_13to17_13), .out_c(matrixC16_13));
processing_element pe16_14(.reset(effective_rst), .clk(clk),  .in_a(a16_13to16_14), .in_b(b15_14to16_14),  .out_a(a16_14to16_15), .out_b(b16_14to17_14), .out_c(matrixC16_14));
processing_element pe16_15(.reset(effective_rst), .clk(clk),  .in_a(a16_14to16_15), .in_b(b15_15to16_15),  .out_a(a16_15to16_16), .out_b(b16_15to17_15), .out_c(matrixC16_15));
processing_element pe16_16(.reset(effective_rst), .clk(clk),  .in_a(a16_15to16_16), .in_b(b15_16to16_16),  .out_a(a16_16to16_17), .out_b(b16_16to17_16), .out_c(matrixC16_16));
processing_element pe16_17(.reset(effective_rst), .clk(clk),  .in_a(a16_16to16_17), .in_b(b15_17to16_17),  .out_a(a16_17to16_18), .out_b(b16_17to17_17), .out_c(matrixC16_17));
processing_element pe16_18(.reset(effective_rst), .clk(clk),  .in_a(a16_17to16_18), .in_b(b15_18to16_18),  .out_a(a16_18to16_19), .out_b(b16_18to17_18), .out_c(matrixC16_18));
processing_element pe16_19(.reset(effective_rst), .clk(clk),  .in_a(a16_18to16_19), .in_b(b15_19to16_19),  .out_a(a16_19to16_20), .out_b(b16_19to17_19), .out_c(matrixC16_19));
processing_element pe16_20(.reset(effective_rst), .clk(clk),  .in_a(a16_19to16_20), .in_b(b15_20to16_20),  .out_a(a16_20to16_21), .out_b(b16_20to17_20), .out_c(matrixC16_20));
processing_element pe16_21(.reset(effective_rst), .clk(clk),  .in_a(a16_20to16_21), .in_b(b15_21to16_21),  .out_a(a16_21to16_22), .out_b(b16_21to17_21), .out_c(matrixC16_21));
processing_element pe16_22(.reset(effective_rst), .clk(clk),  .in_a(a16_21to16_22), .in_b(b15_22to16_22),  .out_a(a16_22to16_23), .out_b(b16_22to17_22), .out_c(matrixC16_22));
processing_element pe16_23(.reset(effective_rst), .clk(clk),  .in_a(a16_22to16_23), .in_b(b15_23to16_23),  .out_a(a16_23to16_24), .out_b(b16_23to17_23), .out_c(matrixC16_23));
processing_element pe16_24(.reset(effective_rst), .clk(clk),  .in_a(a16_23to16_24), .in_b(b15_24to16_24),  .out_a(a16_24to16_25), .out_b(b16_24to17_24), .out_c(matrixC16_24));
processing_element pe16_25(.reset(effective_rst), .clk(clk),  .in_a(a16_24to16_25), .in_b(b15_25to16_25),  .out_a(a16_25to16_26), .out_b(b16_25to17_25), .out_c(matrixC16_25));
processing_element pe16_26(.reset(effective_rst), .clk(clk),  .in_a(a16_25to16_26), .in_b(b15_26to16_26),  .out_a(a16_26to16_27), .out_b(b16_26to17_26), .out_c(matrixC16_26));
processing_element pe16_27(.reset(effective_rst), .clk(clk),  .in_a(a16_26to16_27), .in_b(b15_27to16_27),  .out_a(a16_27to16_28), .out_b(b16_27to17_27), .out_c(matrixC16_27));
processing_element pe16_28(.reset(effective_rst), .clk(clk),  .in_a(a16_27to16_28), .in_b(b15_28to16_28),  .out_a(a16_28to16_29), .out_b(b16_28to17_28), .out_c(matrixC16_28));
processing_element pe16_29(.reset(effective_rst), .clk(clk),  .in_a(a16_28to16_29), .in_b(b15_29to16_29),  .out_a(a16_29to16_30), .out_b(b16_29to17_29), .out_c(matrixC16_29));
processing_element pe16_30(.reset(effective_rst), .clk(clk),  .in_a(a16_29to16_30), .in_b(b15_30to16_30),  .out_a(a16_30to16_31), .out_b(b16_30to17_30), .out_c(matrixC16_30));
processing_element pe16_31(.reset(effective_rst), .clk(clk),  .in_a(a16_30to16_31), .in_b(b15_31to16_31),  .out_a(a16_31to16_32), .out_b(b16_31to17_31), .out_c(matrixC16_31));
processing_element pe17_1(.reset(effective_rst), .clk(clk),  .in_a(a17_0to17_1), .in_b(b16_1to17_1),  .out_a(a17_1to17_2), .out_b(b17_1to18_1), .out_c(matrixC17_1));
processing_element pe17_2(.reset(effective_rst), .clk(clk),  .in_a(a17_1to17_2), .in_b(b16_2to17_2),  .out_a(a17_2to17_3), .out_b(b17_2to18_2), .out_c(matrixC17_2));
processing_element pe17_3(.reset(effective_rst), .clk(clk),  .in_a(a17_2to17_3), .in_b(b16_3to17_3),  .out_a(a17_3to17_4), .out_b(b17_3to18_3), .out_c(matrixC17_3));
processing_element pe17_4(.reset(effective_rst), .clk(clk),  .in_a(a17_3to17_4), .in_b(b16_4to17_4),  .out_a(a17_4to17_5), .out_b(b17_4to18_4), .out_c(matrixC17_4));
processing_element pe17_5(.reset(effective_rst), .clk(clk),  .in_a(a17_4to17_5), .in_b(b16_5to17_5),  .out_a(a17_5to17_6), .out_b(b17_5to18_5), .out_c(matrixC17_5));
processing_element pe17_6(.reset(effective_rst), .clk(clk),  .in_a(a17_5to17_6), .in_b(b16_6to17_6),  .out_a(a17_6to17_7), .out_b(b17_6to18_6), .out_c(matrixC17_6));
processing_element pe17_7(.reset(effective_rst), .clk(clk),  .in_a(a17_6to17_7), .in_b(b16_7to17_7),  .out_a(a17_7to17_8), .out_b(b17_7to18_7), .out_c(matrixC17_7));
processing_element pe17_8(.reset(effective_rst), .clk(clk),  .in_a(a17_7to17_8), .in_b(b16_8to17_8),  .out_a(a17_8to17_9), .out_b(b17_8to18_8), .out_c(matrixC17_8));
processing_element pe17_9(.reset(effective_rst), .clk(clk),  .in_a(a17_8to17_9), .in_b(b16_9to17_9),  .out_a(a17_9to17_10), .out_b(b17_9to18_9), .out_c(matrixC17_9));
processing_element pe17_10(.reset(effective_rst), .clk(clk),  .in_a(a17_9to17_10), .in_b(b16_10to17_10),  .out_a(a17_10to17_11), .out_b(b17_10to18_10), .out_c(matrixC17_10));
processing_element pe17_11(.reset(effective_rst), .clk(clk),  .in_a(a17_10to17_11), .in_b(b16_11to17_11),  .out_a(a17_11to17_12), .out_b(b17_11to18_11), .out_c(matrixC17_11));
processing_element pe17_12(.reset(effective_rst), .clk(clk),  .in_a(a17_11to17_12), .in_b(b16_12to17_12),  .out_a(a17_12to17_13), .out_b(b17_12to18_12), .out_c(matrixC17_12));
processing_element pe17_13(.reset(effective_rst), .clk(clk),  .in_a(a17_12to17_13), .in_b(b16_13to17_13),  .out_a(a17_13to17_14), .out_b(b17_13to18_13), .out_c(matrixC17_13));
processing_element pe17_14(.reset(effective_rst), .clk(clk),  .in_a(a17_13to17_14), .in_b(b16_14to17_14),  .out_a(a17_14to17_15), .out_b(b17_14to18_14), .out_c(matrixC17_14));
processing_element pe17_15(.reset(effective_rst), .clk(clk),  .in_a(a17_14to17_15), .in_b(b16_15to17_15),  .out_a(a17_15to17_16), .out_b(b17_15to18_15), .out_c(matrixC17_15));
processing_element pe17_16(.reset(effective_rst), .clk(clk),  .in_a(a17_15to17_16), .in_b(b16_16to17_16),  .out_a(a17_16to17_17), .out_b(b17_16to18_16), .out_c(matrixC17_16));
processing_element pe17_17(.reset(effective_rst), .clk(clk),  .in_a(a17_16to17_17), .in_b(b16_17to17_17),  .out_a(a17_17to17_18), .out_b(b17_17to18_17), .out_c(matrixC17_17));
processing_element pe17_18(.reset(effective_rst), .clk(clk),  .in_a(a17_17to17_18), .in_b(b16_18to17_18),  .out_a(a17_18to17_19), .out_b(b17_18to18_18), .out_c(matrixC17_18));
processing_element pe17_19(.reset(effective_rst), .clk(clk),  .in_a(a17_18to17_19), .in_b(b16_19to17_19),  .out_a(a17_19to17_20), .out_b(b17_19to18_19), .out_c(matrixC17_19));
processing_element pe17_20(.reset(effective_rst), .clk(clk),  .in_a(a17_19to17_20), .in_b(b16_20to17_20),  .out_a(a17_20to17_21), .out_b(b17_20to18_20), .out_c(matrixC17_20));
processing_element pe17_21(.reset(effective_rst), .clk(clk),  .in_a(a17_20to17_21), .in_b(b16_21to17_21),  .out_a(a17_21to17_22), .out_b(b17_21to18_21), .out_c(matrixC17_21));
processing_element pe17_22(.reset(effective_rst), .clk(clk),  .in_a(a17_21to17_22), .in_b(b16_22to17_22),  .out_a(a17_22to17_23), .out_b(b17_22to18_22), .out_c(matrixC17_22));
processing_element pe17_23(.reset(effective_rst), .clk(clk),  .in_a(a17_22to17_23), .in_b(b16_23to17_23),  .out_a(a17_23to17_24), .out_b(b17_23to18_23), .out_c(matrixC17_23));
processing_element pe17_24(.reset(effective_rst), .clk(clk),  .in_a(a17_23to17_24), .in_b(b16_24to17_24),  .out_a(a17_24to17_25), .out_b(b17_24to18_24), .out_c(matrixC17_24));
processing_element pe17_25(.reset(effective_rst), .clk(clk),  .in_a(a17_24to17_25), .in_b(b16_25to17_25),  .out_a(a17_25to17_26), .out_b(b17_25to18_25), .out_c(matrixC17_25));
processing_element pe17_26(.reset(effective_rst), .clk(clk),  .in_a(a17_25to17_26), .in_b(b16_26to17_26),  .out_a(a17_26to17_27), .out_b(b17_26to18_26), .out_c(matrixC17_26));
processing_element pe17_27(.reset(effective_rst), .clk(clk),  .in_a(a17_26to17_27), .in_b(b16_27to17_27),  .out_a(a17_27to17_28), .out_b(b17_27to18_27), .out_c(matrixC17_27));
processing_element pe17_28(.reset(effective_rst), .clk(clk),  .in_a(a17_27to17_28), .in_b(b16_28to17_28),  .out_a(a17_28to17_29), .out_b(b17_28to18_28), .out_c(matrixC17_28));
processing_element pe17_29(.reset(effective_rst), .clk(clk),  .in_a(a17_28to17_29), .in_b(b16_29to17_29),  .out_a(a17_29to17_30), .out_b(b17_29to18_29), .out_c(matrixC17_29));
processing_element pe17_30(.reset(effective_rst), .clk(clk),  .in_a(a17_29to17_30), .in_b(b16_30to17_30),  .out_a(a17_30to17_31), .out_b(b17_30to18_30), .out_c(matrixC17_30));
processing_element pe17_31(.reset(effective_rst), .clk(clk),  .in_a(a17_30to17_31), .in_b(b16_31to17_31),  .out_a(a17_31to17_32), .out_b(b17_31to18_31), .out_c(matrixC17_31));
processing_element pe18_1(.reset(effective_rst), .clk(clk),  .in_a(a18_0to18_1), .in_b(b17_1to18_1),  .out_a(a18_1to18_2), .out_b(b18_1to19_1), .out_c(matrixC18_1));
processing_element pe18_2(.reset(effective_rst), .clk(clk),  .in_a(a18_1to18_2), .in_b(b17_2to18_2),  .out_a(a18_2to18_3), .out_b(b18_2to19_2), .out_c(matrixC18_2));
processing_element pe18_3(.reset(effective_rst), .clk(clk),  .in_a(a18_2to18_3), .in_b(b17_3to18_3),  .out_a(a18_3to18_4), .out_b(b18_3to19_3), .out_c(matrixC18_3));
processing_element pe18_4(.reset(effective_rst), .clk(clk),  .in_a(a18_3to18_4), .in_b(b17_4to18_4),  .out_a(a18_4to18_5), .out_b(b18_4to19_4), .out_c(matrixC18_4));
processing_element pe18_5(.reset(effective_rst), .clk(clk),  .in_a(a18_4to18_5), .in_b(b17_5to18_5),  .out_a(a18_5to18_6), .out_b(b18_5to19_5), .out_c(matrixC18_5));
processing_element pe18_6(.reset(effective_rst), .clk(clk),  .in_a(a18_5to18_6), .in_b(b17_6to18_6),  .out_a(a18_6to18_7), .out_b(b18_6to19_6), .out_c(matrixC18_6));
processing_element pe18_7(.reset(effective_rst), .clk(clk),  .in_a(a18_6to18_7), .in_b(b17_7to18_7),  .out_a(a18_7to18_8), .out_b(b18_7to19_7), .out_c(matrixC18_7));
processing_element pe18_8(.reset(effective_rst), .clk(clk),  .in_a(a18_7to18_8), .in_b(b17_8to18_8),  .out_a(a18_8to18_9), .out_b(b18_8to19_8), .out_c(matrixC18_8));
processing_element pe18_9(.reset(effective_rst), .clk(clk),  .in_a(a18_8to18_9), .in_b(b17_9to18_9),  .out_a(a18_9to18_10), .out_b(b18_9to19_9), .out_c(matrixC18_9));
processing_element pe18_10(.reset(effective_rst), .clk(clk),  .in_a(a18_9to18_10), .in_b(b17_10to18_10),  .out_a(a18_10to18_11), .out_b(b18_10to19_10), .out_c(matrixC18_10));
processing_element pe18_11(.reset(effective_rst), .clk(clk),  .in_a(a18_10to18_11), .in_b(b17_11to18_11),  .out_a(a18_11to18_12), .out_b(b18_11to19_11), .out_c(matrixC18_11));
processing_element pe18_12(.reset(effective_rst), .clk(clk),  .in_a(a18_11to18_12), .in_b(b17_12to18_12),  .out_a(a18_12to18_13), .out_b(b18_12to19_12), .out_c(matrixC18_12));
processing_element pe18_13(.reset(effective_rst), .clk(clk),  .in_a(a18_12to18_13), .in_b(b17_13to18_13),  .out_a(a18_13to18_14), .out_b(b18_13to19_13), .out_c(matrixC18_13));
processing_element pe18_14(.reset(effective_rst), .clk(clk),  .in_a(a18_13to18_14), .in_b(b17_14to18_14),  .out_a(a18_14to18_15), .out_b(b18_14to19_14), .out_c(matrixC18_14));
processing_element pe18_15(.reset(effective_rst), .clk(clk),  .in_a(a18_14to18_15), .in_b(b17_15to18_15),  .out_a(a18_15to18_16), .out_b(b18_15to19_15), .out_c(matrixC18_15));
processing_element pe18_16(.reset(effective_rst), .clk(clk),  .in_a(a18_15to18_16), .in_b(b17_16to18_16),  .out_a(a18_16to18_17), .out_b(b18_16to19_16), .out_c(matrixC18_16));
processing_element pe18_17(.reset(effective_rst), .clk(clk),  .in_a(a18_16to18_17), .in_b(b17_17to18_17),  .out_a(a18_17to18_18), .out_b(b18_17to19_17), .out_c(matrixC18_17));
processing_element pe18_18(.reset(effective_rst), .clk(clk),  .in_a(a18_17to18_18), .in_b(b17_18to18_18),  .out_a(a18_18to18_19), .out_b(b18_18to19_18), .out_c(matrixC18_18));
processing_element pe18_19(.reset(effective_rst), .clk(clk),  .in_a(a18_18to18_19), .in_b(b17_19to18_19),  .out_a(a18_19to18_20), .out_b(b18_19to19_19), .out_c(matrixC18_19));
processing_element pe18_20(.reset(effective_rst), .clk(clk),  .in_a(a18_19to18_20), .in_b(b17_20to18_20),  .out_a(a18_20to18_21), .out_b(b18_20to19_20), .out_c(matrixC18_20));
processing_element pe18_21(.reset(effective_rst), .clk(clk),  .in_a(a18_20to18_21), .in_b(b17_21to18_21),  .out_a(a18_21to18_22), .out_b(b18_21to19_21), .out_c(matrixC18_21));
processing_element pe18_22(.reset(effective_rst), .clk(clk),  .in_a(a18_21to18_22), .in_b(b17_22to18_22),  .out_a(a18_22to18_23), .out_b(b18_22to19_22), .out_c(matrixC18_22));
processing_element pe18_23(.reset(effective_rst), .clk(clk),  .in_a(a18_22to18_23), .in_b(b17_23to18_23),  .out_a(a18_23to18_24), .out_b(b18_23to19_23), .out_c(matrixC18_23));
processing_element pe18_24(.reset(effective_rst), .clk(clk),  .in_a(a18_23to18_24), .in_b(b17_24to18_24),  .out_a(a18_24to18_25), .out_b(b18_24to19_24), .out_c(matrixC18_24));
processing_element pe18_25(.reset(effective_rst), .clk(clk),  .in_a(a18_24to18_25), .in_b(b17_25to18_25),  .out_a(a18_25to18_26), .out_b(b18_25to19_25), .out_c(matrixC18_25));
processing_element pe18_26(.reset(effective_rst), .clk(clk),  .in_a(a18_25to18_26), .in_b(b17_26to18_26),  .out_a(a18_26to18_27), .out_b(b18_26to19_26), .out_c(matrixC18_26));
processing_element pe18_27(.reset(effective_rst), .clk(clk),  .in_a(a18_26to18_27), .in_b(b17_27to18_27),  .out_a(a18_27to18_28), .out_b(b18_27to19_27), .out_c(matrixC18_27));
processing_element pe18_28(.reset(effective_rst), .clk(clk),  .in_a(a18_27to18_28), .in_b(b17_28to18_28),  .out_a(a18_28to18_29), .out_b(b18_28to19_28), .out_c(matrixC18_28));
processing_element pe18_29(.reset(effective_rst), .clk(clk),  .in_a(a18_28to18_29), .in_b(b17_29to18_29),  .out_a(a18_29to18_30), .out_b(b18_29to19_29), .out_c(matrixC18_29));
processing_element pe18_30(.reset(effective_rst), .clk(clk),  .in_a(a18_29to18_30), .in_b(b17_30to18_30),  .out_a(a18_30to18_31), .out_b(b18_30to19_30), .out_c(matrixC18_30));
processing_element pe18_31(.reset(effective_rst), .clk(clk),  .in_a(a18_30to18_31), .in_b(b17_31to18_31),  .out_a(a18_31to18_32), .out_b(b18_31to19_31), .out_c(matrixC18_31));
processing_element pe19_1(.reset(effective_rst), .clk(clk),  .in_a(a19_0to19_1), .in_b(b18_1to19_1),  .out_a(a19_1to19_2), .out_b(b19_1to20_1), .out_c(matrixC19_1));
processing_element pe19_2(.reset(effective_rst), .clk(clk),  .in_a(a19_1to19_2), .in_b(b18_2to19_2),  .out_a(a19_2to19_3), .out_b(b19_2to20_2), .out_c(matrixC19_2));
processing_element pe19_3(.reset(effective_rst), .clk(clk),  .in_a(a19_2to19_3), .in_b(b18_3to19_3),  .out_a(a19_3to19_4), .out_b(b19_3to20_3), .out_c(matrixC19_3));
processing_element pe19_4(.reset(effective_rst), .clk(clk),  .in_a(a19_3to19_4), .in_b(b18_4to19_4),  .out_a(a19_4to19_5), .out_b(b19_4to20_4), .out_c(matrixC19_4));
processing_element pe19_5(.reset(effective_rst), .clk(clk),  .in_a(a19_4to19_5), .in_b(b18_5to19_5),  .out_a(a19_5to19_6), .out_b(b19_5to20_5), .out_c(matrixC19_5));
processing_element pe19_6(.reset(effective_rst), .clk(clk),  .in_a(a19_5to19_6), .in_b(b18_6to19_6),  .out_a(a19_6to19_7), .out_b(b19_6to20_6), .out_c(matrixC19_6));
processing_element pe19_7(.reset(effective_rst), .clk(clk),  .in_a(a19_6to19_7), .in_b(b18_7to19_7),  .out_a(a19_7to19_8), .out_b(b19_7to20_7), .out_c(matrixC19_7));
processing_element pe19_8(.reset(effective_rst), .clk(clk),  .in_a(a19_7to19_8), .in_b(b18_8to19_8),  .out_a(a19_8to19_9), .out_b(b19_8to20_8), .out_c(matrixC19_8));
processing_element pe19_9(.reset(effective_rst), .clk(clk),  .in_a(a19_8to19_9), .in_b(b18_9to19_9),  .out_a(a19_9to19_10), .out_b(b19_9to20_9), .out_c(matrixC19_9));
processing_element pe19_10(.reset(effective_rst), .clk(clk),  .in_a(a19_9to19_10), .in_b(b18_10to19_10),  .out_a(a19_10to19_11), .out_b(b19_10to20_10), .out_c(matrixC19_10));
processing_element pe19_11(.reset(effective_rst), .clk(clk),  .in_a(a19_10to19_11), .in_b(b18_11to19_11),  .out_a(a19_11to19_12), .out_b(b19_11to20_11), .out_c(matrixC19_11));
processing_element pe19_12(.reset(effective_rst), .clk(clk),  .in_a(a19_11to19_12), .in_b(b18_12to19_12),  .out_a(a19_12to19_13), .out_b(b19_12to20_12), .out_c(matrixC19_12));
processing_element pe19_13(.reset(effective_rst), .clk(clk),  .in_a(a19_12to19_13), .in_b(b18_13to19_13),  .out_a(a19_13to19_14), .out_b(b19_13to20_13), .out_c(matrixC19_13));
processing_element pe19_14(.reset(effective_rst), .clk(clk),  .in_a(a19_13to19_14), .in_b(b18_14to19_14),  .out_a(a19_14to19_15), .out_b(b19_14to20_14), .out_c(matrixC19_14));
processing_element pe19_15(.reset(effective_rst), .clk(clk),  .in_a(a19_14to19_15), .in_b(b18_15to19_15),  .out_a(a19_15to19_16), .out_b(b19_15to20_15), .out_c(matrixC19_15));
processing_element pe19_16(.reset(effective_rst), .clk(clk),  .in_a(a19_15to19_16), .in_b(b18_16to19_16),  .out_a(a19_16to19_17), .out_b(b19_16to20_16), .out_c(matrixC19_16));
processing_element pe19_17(.reset(effective_rst), .clk(clk),  .in_a(a19_16to19_17), .in_b(b18_17to19_17),  .out_a(a19_17to19_18), .out_b(b19_17to20_17), .out_c(matrixC19_17));
processing_element pe19_18(.reset(effective_rst), .clk(clk),  .in_a(a19_17to19_18), .in_b(b18_18to19_18),  .out_a(a19_18to19_19), .out_b(b19_18to20_18), .out_c(matrixC19_18));
processing_element pe19_19(.reset(effective_rst), .clk(clk),  .in_a(a19_18to19_19), .in_b(b18_19to19_19),  .out_a(a19_19to19_20), .out_b(b19_19to20_19), .out_c(matrixC19_19));
processing_element pe19_20(.reset(effective_rst), .clk(clk),  .in_a(a19_19to19_20), .in_b(b18_20to19_20),  .out_a(a19_20to19_21), .out_b(b19_20to20_20), .out_c(matrixC19_20));
processing_element pe19_21(.reset(effective_rst), .clk(clk),  .in_a(a19_20to19_21), .in_b(b18_21to19_21),  .out_a(a19_21to19_22), .out_b(b19_21to20_21), .out_c(matrixC19_21));
processing_element pe19_22(.reset(effective_rst), .clk(clk),  .in_a(a19_21to19_22), .in_b(b18_22to19_22),  .out_a(a19_22to19_23), .out_b(b19_22to20_22), .out_c(matrixC19_22));
processing_element pe19_23(.reset(effective_rst), .clk(clk),  .in_a(a19_22to19_23), .in_b(b18_23to19_23),  .out_a(a19_23to19_24), .out_b(b19_23to20_23), .out_c(matrixC19_23));
processing_element pe19_24(.reset(effective_rst), .clk(clk),  .in_a(a19_23to19_24), .in_b(b18_24to19_24),  .out_a(a19_24to19_25), .out_b(b19_24to20_24), .out_c(matrixC19_24));
processing_element pe19_25(.reset(effective_rst), .clk(clk),  .in_a(a19_24to19_25), .in_b(b18_25to19_25),  .out_a(a19_25to19_26), .out_b(b19_25to20_25), .out_c(matrixC19_25));
processing_element pe19_26(.reset(effective_rst), .clk(clk),  .in_a(a19_25to19_26), .in_b(b18_26to19_26),  .out_a(a19_26to19_27), .out_b(b19_26to20_26), .out_c(matrixC19_26));
processing_element pe19_27(.reset(effective_rst), .clk(clk),  .in_a(a19_26to19_27), .in_b(b18_27to19_27),  .out_a(a19_27to19_28), .out_b(b19_27to20_27), .out_c(matrixC19_27));
processing_element pe19_28(.reset(effective_rst), .clk(clk),  .in_a(a19_27to19_28), .in_b(b18_28to19_28),  .out_a(a19_28to19_29), .out_b(b19_28to20_28), .out_c(matrixC19_28));
processing_element pe19_29(.reset(effective_rst), .clk(clk),  .in_a(a19_28to19_29), .in_b(b18_29to19_29),  .out_a(a19_29to19_30), .out_b(b19_29to20_29), .out_c(matrixC19_29));
processing_element pe19_30(.reset(effective_rst), .clk(clk),  .in_a(a19_29to19_30), .in_b(b18_30to19_30),  .out_a(a19_30to19_31), .out_b(b19_30to20_30), .out_c(matrixC19_30));
processing_element pe19_31(.reset(effective_rst), .clk(clk),  .in_a(a19_30to19_31), .in_b(b18_31to19_31),  .out_a(a19_31to19_32), .out_b(b19_31to20_31), .out_c(matrixC19_31));
processing_element pe20_1(.reset(effective_rst), .clk(clk),  .in_a(a20_0to20_1), .in_b(b19_1to20_1),  .out_a(a20_1to20_2), .out_b(b20_1to21_1), .out_c(matrixC20_1));
processing_element pe20_2(.reset(effective_rst), .clk(clk),  .in_a(a20_1to20_2), .in_b(b19_2to20_2),  .out_a(a20_2to20_3), .out_b(b20_2to21_2), .out_c(matrixC20_2));
processing_element pe20_3(.reset(effective_rst), .clk(clk),  .in_a(a20_2to20_3), .in_b(b19_3to20_3),  .out_a(a20_3to20_4), .out_b(b20_3to21_3), .out_c(matrixC20_3));
processing_element pe20_4(.reset(effective_rst), .clk(clk),  .in_a(a20_3to20_4), .in_b(b19_4to20_4),  .out_a(a20_4to20_5), .out_b(b20_4to21_4), .out_c(matrixC20_4));
processing_element pe20_5(.reset(effective_rst), .clk(clk),  .in_a(a20_4to20_5), .in_b(b19_5to20_5),  .out_a(a20_5to20_6), .out_b(b20_5to21_5), .out_c(matrixC20_5));
processing_element pe20_6(.reset(effective_rst), .clk(clk),  .in_a(a20_5to20_6), .in_b(b19_6to20_6),  .out_a(a20_6to20_7), .out_b(b20_6to21_6), .out_c(matrixC20_6));
processing_element pe20_7(.reset(effective_rst), .clk(clk),  .in_a(a20_6to20_7), .in_b(b19_7to20_7),  .out_a(a20_7to20_8), .out_b(b20_7to21_7), .out_c(matrixC20_7));
processing_element pe20_8(.reset(effective_rst), .clk(clk),  .in_a(a20_7to20_8), .in_b(b19_8to20_8),  .out_a(a20_8to20_9), .out_b(b20_8to21_8), .out_c(matrixC20_8));
processing_element pe20_9(.reset(effective_rst), .clk(clk),  .in_a(a20_8to20_9), .in_b(b19_9to20_9),  .out_a(a20_9to20_10), .out_b(b20_9to21_9), .out_c(matrixC20_9));
processing_element pe20_10(.reset(effective_rst), .clk(clk),  .in_a(a20_9to20_10), .in_b(b19_10to20_10),  .out_a(a20_10to20_11), .out_b(b20_10to21_10), .out_c(matrixC20_10));
processing_element pe20_11(.reset(effective_rst), .clk(clk),  .in_a(a20_10to20_11), .in_b(b19_11to20_11),  .out_a(a20_11to20_12), .out_b(b20_11to21_11), .out_c(matrixC20_11));
processing_element pe20_12(.reset(effective_rst), .clk(clk),  .in_a(a20_11to20_12), .in_b(b19_12to20_12),  .out_a(a20_12to20_13), .out_b(b20_12to21_12), .out_c(matrixC20_12));
processing_element pe20_13(.reset(effective_rst), .clk(clk),  .in_a(a20_12to20_13), .in_b(b19_13to20_13),  .out_a(a20_13to20_14), .out_b(b20_13to21_13), .out_c(matrixC20_13));
processing_element pe20_14(.reset(effective_rst), .clk(clk),  .in_a(a20_13to20_14), .in_b(b19_14to20_14),  .out_a(a20_14to20_15), .out_b(b20_14to21_14), .out_c(matrixC20_14));
processing_element pe20_15(.reset(effective_rst), .clk(clk),  .in_a(a20_14to20_15), .in_b(b19_15to20_15),  .out_a(a20_15to20_16), .out_b(b20_15to21_15), .out_c(matrixC20_15));
processing_element pe20_16(.reset(effective_rst), .clk(clk),  .in_a(a20_15to20_16), .in_b(b19_16to20_16),  .out_a(a20_16to20_17), .out_b(b20_16to21_16), .out_c(matrixC20_16));
processing_element pe20_17(.reset(effective_rst), .clk(clk),  .in_a(a20_16to20_17), .in_b(b19_17to20_17),  .out_a(a20_17to20_18), .out_b(b20_17to21_17), .out_c(matrixC20_17));
processing_element pe20_18(.reset(effective_rst), .clk(clk),  .in_a(a20_17to20_18), .in_b(b19_18to20_18),  .out_a(a20_18to20_19), .out_b(b20_18to21_18), .out_c(matrixC20_18));
processing_element pe20_19(.reset(effective_rst), .clk(clk),  .in_a(a20_18to20_19), .in_b(b19_19to20_19),  .out_a(a20_19to20_20), .out_b(b20_19to21_19), .out_c(matrixC20_19));
processing_element pe20_20(.reset(effective_rst), .clk(clk),  .in_a(a20_19to20_20), .in_b(b19_20to20_20),  .out_a(a20_20to20_21), .out_b(b20_20to21_20), .out_c(matrixC20_20));
processing_element pe20_21(.reset(effective_rst), .clk(clk),  .in_a(a20_20to20_21), .in_b(b19_21to20_21),  .out_a(a20_21to20_22), .out_b(b20_21to21_21), .out_c(matrixC20_21));
processing_element pe20_22(.reset(effective_rst), .clk(clk),  .in_a(a20_21to20_22), .in_b(b19_22to20_22),  .out_a(a20_22to20_23), .out_b(b20_22to21_22), .out_c(matrixC20_22));
processing_element pe20_23(.reset(effective_rst), .clk(clk),  .in_a(a20_22to20_23), .in_b(b19_23to20_23),  .out_a(a20_23to20_24), .out_b(b20_23to21_23), .out_c(matrixC20_23));
processing_element pe20_24(.reset(effective_rst), .clk(clk),  .in_a(a20_23to20_24), .in_b(b19_24to20_24),  .out_a(a20_24to20_25), .out_b(b20_24to21_24), .out_c(matrixC20_24));
processing_element pe20_25(.reset(effective_rst), .clk(clk),  .in_a(a20_24to20_25), .in_b(b19_25to20_25),  .out_a(a20_25to20_26), .out_b(b20_25to21_25), .out_c(matrixC20_25));
processing_element pe20_26(.reset(effective_rst), .clk(clk),  .in_a(a20_25to20_26), .in_b(b19_26to20_26),  .out_a(a20_26to20_27), .out_b(b20_26to21_26), .out_c(matrixC20_26));
processing_element pe20_27(.reset(effective_rst), .clk(clk),  .in_a(a20_26to20_27), .in_b(b19_27to20_27),  .out_a(a20_27to20_28), .out_b(b20_27to21_27), .out_c(matrixC20_27));
processing_element pe20_28(.reset(effective_rst), .clk(clk),  .in_a(a20_27to20_28), .in_b(b19_28to20_28),  .out_a(a20_28to20_29), .out_b(b20_28to21_28), .out_c(matrixC20_28));
processing_element pe20_29(.reset(effective_rst), .clk(clk),  .in_a(a20_28to20_29), .in_b(b19_29to20_29),  .out_a(a20_29to20_30), .out_b(b20_29to21_29), .out_c(matrixC20_29));
processing_element pe20_30(.reset(effective_rst), .clk(clk),  .in_a(a20_29to20_30), .in_b(b19_30to20_30),  .out_a(a20_30to20_31), .out_b(b20_30to21_30), .out_c(matrixC20_30));
processing_element pe20_31(.reset(effective_rst), .clk(clk),  .in_a(a20_30to20_31), .in_b(b19_31to20_31),  .out_a(a20_31to20_32), .out_b(b20_31to21_31), .out_c(matrixC20_31));
processing_element pe21_1(.reset(effective_rst), .clk(clk),  .in_a(a21_0to21_1), .in_b(b20_1to21_1),  .out_a(a21_1to21_2), .out_b(b21_1to22_1), .out_c(matrixC21_1));
processing_element pe21_2(.reset(effective_rst), .clk(clk),  .in_a(a21_1to21_2), .in_b(b20_2to21_2),  .out_a(a21_2to21_3), .out_b(b21_2to22_2), .out_c(matrixC21_2));
processing_element pe21_3(.reset(effective_rst), .clk(clk),  .in_a(a21_2to21_3), .in_b(b20_3to21_3),  .out_a(a21_3to21_4), .out_b(b21_3to22_3), .out_c(matrixC21_3));
processing_element pe21_4(.reset(effective_rst), .clk(clk),  .in_a(a21_3to21_4), .in_b(b20_4to21_4),  .out_a(a21_4to21_5), .out_b(b21_4to22_4), .out_c(matrixC21_4));
processing_element pe21_5(.reset(effective_rst), .clk(clk),  .in_a(a21_4to21_5), .in_b(b20_5to21_5),  .out_a(a21_5to21_6), .out_b(b21_5to22_5), .out_c(matrixC21_5));
processing_element pe21_6(.reset(effective_rst), .clk(clk),  .in_a(a21_5to21_6), .in_b(b20_6to21_6),  .out_a(a21_6to21_7), .out_b(b21_6to22_6), .out_c(matrixC21_6));
processing_element pe21_7(.reset(effective_rst), .clk(clk),  .in_a(a21_6to21_7), .in_b(b20_7to21_7),  .out_a(a21_7to21_8), .out_b(b21_7to22_7), .out_c(matrixC21_7));
processing_element pe21_8(.reset(effective_rst), .clk(clk),  .in_a(a21_7to21_8), .in_b(b20_8to21_8),  .out_a(a21_8to21_9), .out_b(b21_8to22_8), .out_c(matrixC21_8));
processing_element pe21_9(.reset(effective_rst), .clk(clk),  .in_a(a21_8to21_9), .in_b(b20_9to21_9),  .out_a(a21_9to21_10), .out_b(b21_9to22_9), .out_c(matrixC21_9));
processing_element pe21_10(.reset(effective_rst), .clk(clk),  .in_a(a21_9to21_10), .in_b(b20_10to21_10),  .out_a(a21_10to21_11), .out_b(b21_10to22_10), .out_c(matrixC21_10));
processing_element pe21_11(.reset(effective_rst), .clk(clk),  .in_a(a21_10to21_11), .in_b(b20_11to21_11),  .out_a(a21_11to21_12), .out_b(b21_11to22_11), .out_c(matrixC21_11));
processing_element pe21_12(.reset(effective_rst), .clk(clk),  .in_a(a21_11to21_12), .in_b(b20_12to21_12),  .out_a(a21_12to21_13), .out_b(b21_12to22_12), .out_c(matrixC21_12));
processing_element pe21_13(.reset(effective_rst), .clk(clk),  .in_a(a21_12to21_13), .in_b(b20_13to21_13),  .out_a(a21_13to21_14), .out_b(b21_13to22_13), .out_c(matrixC21_13));
processing_element pe21_14(.reset(effective_rst), .clk(clk),  .in_a(a21_13to21_14), .in_b(b20_14to21_14),  .out_a(a21_14to21_15), .out_b(b21_14to22_14), .out_c(matrixC21_14));
processing_element pe21_15(.reset(effective_rst), .clk(clk),  .in_a(a21_14to21_15), .in_b(b20_15to21_15),  .out_a(a21_15to21_16), .out_b(b21_15to22_15), .out_c(matrixC21_15));
processing_element pe21_16(.reset(effective_rst), .clk(clk),  .in_a(a21_15to21_16), .in_b(b20_16to21_16),  .out_a(a21_16to21_17), .out_b(b21_16to22_16), .out_c(matrixC21_16));
processing_element pe21_17(.reset(effective_rst), .clk(clk),  .in_a(a21_16to21_17), .in_b(b20_17to21_17),  .out_a(a21_17to21_18), .out_b(b21_17to22_17), .out_c(matrixC21_17));
processing_element pe21_18(.reset(effective_rst), .clk(clk),  .in_a(a21_17to21_18), .in_b(b20_18to21_18),  .out_a(a21_18to21_19), .out_b(b21_18to22_18), .out_c(matrixC21_18));
processing_element pe21_19(.reset(effective_rst), .clk(clk),  .in_a(a21_18to21_19), .in_b(b20_19to21_19),  .out_a(a21_19to21_20), .out_b(b21_19to22_19), .out_c(matrixC21_19));
processing_element pe21_20(.reset(effective_rst), .clk(clk),  .in_a(a21_19to21_20), .in_b(b20_20to21_20),  .out_a(a21_20to21_21), .out_b(b21_20to22_20), .out_c(matrixC21_20));
processing_element pe21_21(.reset(effective_rst), .clk(clk),  .in_a(a21_20to21_21), .in_b(b20_21to21_21),  .out_a(a21_21to21_22), .out_b(b21_21to22_21), .out_c(matrixC21_21));
processing_element pe21_22(.reset(effective_rst), .clk(clk),  .in_a(a21_21to21_22), .in_b(b20_22to21_22),  .out_a(a21_22to21_23), .out_b(b21_22to22_22), .out_c(matrixC21_22));
processing_element pe21_23(.reset(effective_rst), .clk(clk),  .in_a(a21_22to21_23), .in_b(b20_23to21_23),  .out_a(a21_23to21_24), .out_b(b21_23to22_23), .out_c(matrixC21_23));
processing_element pe21_24(.reset(effective_rst), .clk(clk),  .in_a(a21_23to21_24), .in_b(b20_24to21_24),  .out_a(a21_24to21_25), .out_b(b21_24to22_24), .out_c(matrixC21_24));
processing_element pe21_25(.reset(effective_rst), .clk(clk),  .in_a(a21_24to21_25), .in_b(b20_25to21_25),  .out_a(a21_25to21_26), .out_b(b21_25to22_25), .out_c(matrixC21_25));
processing_element pe21_26(.reset(effective_rst), .clk(clk),  .in_a(a21_25to21_26), .in_b(b20_26to21_26),  .out_a(a21_26to21_27), .out_b(b21_26to22_26), .out_c(matrixC21_26));
processing_element pe21_27(.reset(effective_rst), .clk(clk),  .in_a(a21_26to21_27), .in_b(b20_27to21_27),  .out_a(a21_27to21_28), .out_b(b21_27to22_27), .out_c(matrixC21_27));
processing_element pe21_28(.reset(effective_rst), .clk(clk),  .in_a(a21_27to21_28), .in_b(b20_28to21_28),  .out_a(a21_28to21_29), .out_b(b21_28to22_28), .out_c(matrixC21_28));
processing_element pe21_29(.reset(effective_rst), .clk(clk),  .in_a(a21_28to21_29), .in_b(b20_29to21_29),  .out_a(a21_29to21_30), .out_b(b21_29to22_29), .out_c(matrixC21_29));
processing_element pe21_30(.reset(effective_rst), .clk(clk),  .in_a(a21_29to21_30), .in_b(b20_30to21_30),  .out_a(a21_30to21_31), .out_b(b21_30to22_30), .out_c(matrixC21_30));
processing_element pe21_31(.reset(effective_rst), .clk(clk),  .in_a(a21_30to21_31), .in_b(b20_31to21_31),  .out_a(a21_31to21_32), .out_b(b21_31to22_31), .out_c(matrixC21_31));
processing_element pe22_1(.reset(effective_rst), .clk(clk),  .in_a(a22_0to22_1), .in_b(b21_1to22_1),  .out_a(a22_1to22_2), .out_b(b22_1to23_1), .out_c(matrixC22_1));
processing_element pe22_2(.reset(effective_rst), .clk(clk),  .in_a(a22_1to22_2), .in_b(b21_2to22_2),  .out_a(a22_2to22_3), .out_b(b22_2to23_2), .out_c(matrixC22_2));
processing_element pe22_3(.reset(effective_rst), .clk(clk),  .in_a(a22_2to22_3), .in_b(b21_3to22_3),  .out_a(a22_3to22_4), .out_b(b22_3to23_3), .out_c(matrixC22_3));
processing_element pe22_4(.reset(effective_rst), .clk(clk),  .in_a(a22_3to22_4), .in_b(b21_4to22_4),  .out_a(a22_4to22_5), .out_b(b22_4to23_4), .out_c(matrixC22_4));
processing_element pe22_5(.reset(effective_rst), .clk(clk),  .in_a(a22_4to22_5), .in_b(b21_5to22_5),  .out_a(a22_5to22_6), .out_b(b22_5to23_5), .out_c(matrixC22_5));
processing_element pe22_6(.reset(effective_rst), .clk(clk),  .in_a(a22_5to22_6), .in_b(b21_6to22_6),  .out_a(a22_6to22_7), .out_b(b22_6to23_6), .out_c(matrixC22_6));
processing_element pe22_7(.reset(effective_rst), .clk(clk),  .in_a(a22_6to22_7), .in_b(b21_7to22_7),  .out_a(a22_7to22_8), .out_b(b22_7to23_7), .out_c(matrixC22_7));
processing_element pe22_8(.reset(effective_rst), .clk(clk),  .in_a(a22_7to22_8), .in_b(b21_8to22_8),  .out_a(a22_8to22_9), .out_b(b22_8to23_8), .out_c(matrixC22_8));
processing_element pe22_9(.reset(effective_rst), .clk(clk),  .in_a(a22_8to22_9), .in_b(b21_9to22_9),  .out_a(a22_9to22_10), .out_b(b22_9to23_9), .out_c(matrixC22_9));
processing_element pe22_10(.reset(effective_rst), .clk(clk),  .in_a(a22_9to22_10), .in_b(b21_10to22_10),  .out_a(a22_10to22_11), .out_b(b22_10to23_10), .out_c(matrixC22_10));
processing_element pe22_11(.reset(effective_rst), .clk(clk),  .in_a(a22_10to22_11), .in_b(b21_11to22_11),  .out_a(a22_11to22_12), .out_b(b22_11to23_11), .out_c(matrixC22_11));
processing_element pe22_12(.reset(effective_rst), .clk(clk),  .in_a(a22_11to22_12), .in_b(b21_12to22_12),  .out_a(a22_12to22_13), .out_b(b22_12to23_12), .out_c(matrixC22_12));
processing_element pe22_13(.reset(effective_rst), .clk(clk),  .in_a(a22_12to22_13), .in_b(b21_13to22_13),  .out_a(a22_13to22_14), .out_b(b22_13to23_13), .out_c(matrixC22_13));
processing_element pe22_14(.reset(effective_rst), .clk(clk),  .in_a(a22_13to22_14), .in_b(b21_14to22_14),  .out_a(a22_14to22_15), .out_b(b22_14to23_14), .out_c(matrixC22_14));
processing_element pe22_15(.reset(effective_rst), .clk(clk),  .in_a(a22_14to22_15), .in_b(b21_15to22_15),  .out_a(a22_15to22_16), .out_b(b22_15to23_15), .out_c(matrixC22_15));
processing_element pe22_16(.reset(effective_rst), .clk(clk),  .in_a(a22_15to22_16), .in_b(b21_16to22_16),  .out_a(a22_16to22_17), .out_b(b22_16to23_16), .out_c(matrixC22_16));
processing_element pe22_17(.reset(effective_rst), .clk(clk),  .in_a(a22_16to22_17), .in_b(b21_17to22_17),  .out_a(a22_17to22_18), .out_b(b22_17to23_17), .out_c(matrixC22_17));
processing_element pe22_18(.reset(effective_rst), .clk(clk),  .in_a(a22_17to22_18), .in_b(b21_18to22_18),  .out_a(a22_18to22_19), .out_b(b22_18to23_18), .out_c(matrixC22_18));
processing_element pe22_19(.reset(effective_rst), .clk(clk),  .in_a(a22_18to22_19), .in_b(b21_19to22_19),  .out_a(a22_19to22_20), .out_b(b22_19to23_19), .out_c(matrixC22_19));
processing_element pe22_20(.reset(effective_rst), .clk(clk),  .in_a(a22_19to22_20), .in_b(b21_20to22_20),  .out_a(a22_20to22_21), .out_b(b22_20to23_20), .out_c(matrixC22_20));
processing_element pe22_21(.reset(effective_rst), .clk(clk),  .in_a(a22_20to22_21), .in_b(b21_21to22_21),  .out_a(a22_21to22_22), .out_b(b22_21to23_21), .out_c(matrixC22_21));
processing_element pe22_22(.reset(effective_rst), .clk(clk),  .in_a(a22_21to22_22), .in_b(b21_22to22_22),  .out_a(a22_22to22_23), .out_b(b22_22to23_22), .out_c(matrixC22_22));
processing_element pe22_23(.reset(effective_rst), .clk(clk),  .in_a(a22_22to22_23), .in_b(b21_23to22_23),  .out_a(a22_23to22_24), .out_b(b22_23to23_23), .out_c(matrixC22_23));
processing_element pe22_24(.reset(effective_rst), .clk(clk),  .in_a(a22_23to22_24), .in_b(b21_24to22_24),  .out_a(a22_24to22_25), .out_b(b22_24to23_24), .out_c(matrixC22_24));
processing_element pe22_25(.reset(effective_rst), .clk(clk),  .in_a(a22_24to22_25), .in_b(b21_25to22_25),  .out_a(a22_25to22_26), .out_b(b22_25to23_25), .out_c(matrixC22_25));
processing_element pe22_26(.reset(effective_rst), .clk(clk),  .in_a(a22_25to22_26), .in_b(b21_26to22_26),  .out_a(a22_26to22_27), .out_b(b22_26to23_26), .out_c(matrixC22_26));
processing_element pe22_27(.reset(effective_rst), .clk(clk),  .in_a(a22_26to22_27), .in_b(b21_27to22_27),  .out_a(a22_27to22_28), .out_b(b22_27to23_27), .out_c(matrixC22_27));
processing_element pe22_28(.reset(effective_rst), .clk(clk),  .in_a(a22_27to22_28), .in_b(b21_28to22_28),  .out_a(a22_28to22_29), .out_b(b22_28to23_28), .out_c(matrixC22_28));
processing_element pe22_29(.reset(effective_rst), .clk(clk),  .in_a(a22_28to22_29), .in_b(b21_29to22_29),  .out_a(a22_29to22_30), .out_b(b22_29to23_29), .out_c(matrixC22_29));
processing_element pe22_30(.reset(effective_rst), .clk(clk),  .in_a(a22_29to22_30), .in_b(b21_30to22_30),  .out_a(a22_30to22_31), .out_b(b22_30to23_30), .out_c(matrixC22_30));
processing_element pe22_31(.reset(effective_rst), .clk(clk),  .in_a(a22_30to22_31), .in_b(b21_31to22_31),  .out_a(a22_31to22_32), .out_b(b22_31to23_31), .out_c(matrixC22_31));
processing_element pe23_1(.reset(effective_rst), .clk(clk),  .in_a(a23_0to23_1), .in_b(b22_1to23_1),  .out_a(a23_1to23_2), .out_b(b23_1to24_1), .out_c(matrixC23_1));
processing_element pe23_2(.reset(effective_rst), .clk(clk),  .in_a(a23_1to23_2), .in_b(b22_2to23_2),  .out_a(a23_2to23_3), .out_b(b23_2to24_2), .out_c(matrixC23_2));
processing_element pe23_3(.reset(effective_rst), .clk(clk),  .in_a(a23_2to23_3), .in_b(b22_3to23_3),  .out_a(a23_3to23_4), .out_b(b23_3to24_3), .out_c(matrixC23_3));
processing_element pe23_4(.reset(effective_rst), .clk(clk),  .in_a(a23_3to23_4), .in_b(b22_4to23_4),  .out_a(a23_4to23_5), .out_b(b23_4to24_4), .out_c(matrixC23_4));
processing_element pe23_5(.reset(effective_rst), .clk(clk),  .in_a(a23_4to23_5), .in_b(b22_5to23_5),  .out_a(a23_5to23_6), .out_b(b23_5to24_5), .out_c(matrixC23_5));
processing_element pe23_6(.reset(effective_rst), .clk(clk),  .in_a(a23_5to23_6), .in_b(b22_6to23_6),  .out_a(a23_6to23_7), .out_b(b23_6to24_6), .out_c(matrixC23_6));
processing_element pe23_7(.reset(effective_rst), .clk(clk),  .in_a(a23_6to23_7), .in_b(b22_7to23_7),  .out_a(a23_7to23_8), .out_b(b23_7to24_7), .out_c(matrixC23_7));
processing_element pe23_8(.reset(effective_rst), .clk(clk),  .in_a(a23_7to23_8), .in_b(b22_8to23_8),  .out_a(a23_8to23_9), .out_b(b23_8to24_8), .out_c(matrixC23_8));
processing_element pe23_9(.reset(effective_rst), .clk(clk),  .in_a(a23_8to23_9), .in_b(b22_9to23_9),  .out_a(a23_9to23_10), .out_b(b23_9to24_9), .out_c(matrixC23_9));
processing_element pe23_10(.reset(effective_rst), .clk(clk),  .in_a(a23_9to23_10), .in_b(b22_10to23_10),  .out_a(a23_10to23_11), .out_b(b23_10to24_10), .out_c(matrixC23_10));
processing_element pe23_11(.reset(effective_rst), .clk(clk),  .in_a(a23_10to23_11), .in_b(b22_11to23_11),  .out_a(a23_11to23_12), .out_b(b23_11to24_11), .out_c(matrixC23_11));
processing_element pe23_12(.reset(effective_rst), .clk(clk),  .in_a(a23_11to23_12), .in_b(b22_12to23_12),  .out_a(a23_12to23_13), .out_b(b23_12to24_12), .out_c(matrixC23_12));
processing_element pe23_13(.reset(effective_rst), .clk(clk),  .in_a(a23_12to23_13), .in_b(b22_13to23_13),  .out_a(a23_13to23_14), .out_b(b23_13to24_13), .out_c(matrixC23_13));
processing_element pe23_14(.reset(effective_rst), .clk(clk),  .in_a(a23_13to23_14), .in_b(b22_14to23_14),  .out_a(a23_14to23_15), .out_b(b23_14to24_14), .out_c(matrixC23_14));
processing_element pe23_15(.reset(effective_rst), .clk(clk),  .in_a(a23_14to23_15), .in_b(b22_15to23_15),  .out_a(a23_15to23_16), .out_b(b23_15to24_15), .out_c(matrixC23_15));
processing_element pe23_16(.reset(effective_rst), .clk(clk),  .in_a(a23_15to23_16), .in_b(b22_16to23_16),  .out_a(a23_16to23_17), .out_b(b23_16to24_16), .out_c(matrixC23_16));
processing_element pe23_17(.reset(effective_rst), .clk(clk),  .in_a(a23_16to23_17), .in_b(b22_17to23_17),  .out_a(a23_17to23_18), .out_b(b23_17to24_17), .out_c(matrixC23_17));
processing_element pe23_18(.reset(effective_rst), .clk(clk),  .in_a(a23_17to23_18), .in_b(b22_18to23_18),  .out_a(a23_18to23_19), .out_b(b23_18to24_18), .out_c(matrixC23_18));
processing_element pe23_19(.reset(effective_rst), .clk(clk),  .in_a(a23_18to23_19), .in_b(b22_19to23_19),  .out_a(a23_19to23_20), .out_b(b23_19to24_19), .out_c(matrixC23_19));
processing_element pe23_20(.reset(effective_rst), .clk(clk),  .in_a(a23_19to23_20), .in_b(b22_20to23_20),  .out_a(a23_20to23_21), .out_b(b23_20to24_20), .out_c(matrixC23_20));
processing_element pe23_21(.reset(effective_rst), .clk(clk),  .in_a(a23_20to23_21), .in_b(b22_21to23_21),  .out_a(a23_21to23_22), .out_b(b23_21to24_21), .out_c(matrixC23_21));
processing_element pe23_22(.reset(effective_rst), .clk(clk),  .in_a(a23_21to23_22), .in_b(b22_22to23_22),  .out_a(a23_22to23_23), .out_b(b23_22to24_22), .out_c(matrixC23_22));
processing_element pe23_23(.reset(effective_rst), .clk(clk),  .in_a(a23_22to23_23), .in_b(b22_23to23_23),  .out_a(a23_23to23_24), .out_b(b23_23to24_23), .out_c(matrixC23_23));
processing_element pe23_24(.reset(effective_rst), .clk(clk),  .in_a(a23_23to23_24), .in_b(b22_24to23_24),  .out_a(a23_24to23_25), .out_b(b23_24to24_24), .out_c(matrixC23_24));
processing_element pe23_25(.reset(effective_rst), .clk(clk),  .in_a(a23_24to23_25), .in_b(b22_25to23_25),  .out_a(a23_25to23_26), .out_b(b23_25to24_25), .out_c(matrixC23_25));
processing_element pe23_26(.reset(effective_rst), .clk(clk),  .in_a(a23_25to23_26), .in_b(b22_26to23_26),  .out_a(a23_26to23_27), .out_b(b23_26to24_26), .out_c(matrixC23_26));
processing_element pe23_27(.reset(effective_rst), .clk(clk),  .in_a(a23_26to23_27), .in_b(b22_27to23_27),  .out_a(a23_27to23_28), .out_b(b23_27to24_27), .out_c(matrixC23_27));
processing_element pe23_28(.reset(effective_rst), .clk(clk),  .in_a(a23_27to23_28), .in_b(b22_28to23_28),  .out_a(a23_28to23_29), .out_b(b23_28to24_28), .out_c(matrixC23_28));
processing_element pe23_29(.reset(effective_rst), .clk(clk),  .in_a(a23_28to23_29), .in_b(b22_29to23_29),  .out_a(a23_29to23_30), .out_b(b23_29to24_29), .out_c(matrixC23_29));
processing_element pe23_30(.reset(effective_rst), .clk(clk),  .in_a(a23_29to23_30), .in_b(b22_30to23_30),  .out_a(a23_30to23_31), .out_b(b23_30to24_30), .out_c(matrixC23_30));
processing_element pe23_31(.reset(effective_rst), .clk(clk),  .in_a(a23_30to23_31), .in_b(b22_31to23_31),  .out_a(a23_31to23_32), .out_b(b23_31to24_31), .out_c(matrixC23_31));
processing_element pe24_1(.reset(effective_rst), .clk(clk),  .in_a(a24_0to24_1), .in_b(b23_1to24_1),  .out_a(a24_1to24_2), .out_b(b24_1to25_1), .out_c(matrixC24_1));
processing_element pe24_2(.reset(effective_rst), .clk(clk),  .in_a(a24_1to24_2), .in_b(b23_2to24_2),  .out_a(a24_2to24_3), .out_b(b24_2to25_2), .out_c(matrixC24_2));
processing_element pe24_3(.reset(effective_rst), .clk(clk),  .in_a(a24_2to24_3), .in_b(b23_3to24_3),  .out_a(a24_3to24_4), .out_b(b24_3to25_3), .out_c(matrixC24_3));
processing_element pe24_4(.reset(effective_rst), .clk(clk),  .in_a(a24_3to24_4), .in_b(b23_4to24_4),  .out_a(a24_4to24_5), .out_b(b24_4to25_4), .out_c(matrixC24_4));
processing_element pe24_5(.reset(effective_rst), .clk(clk),  .in_a(a24_4to24_5), .in_b(b23_5to24_5),  .out_a(a24_5to24_6), .out_b(b24_5to25_5), .out_c(matrixC24_5));
processing_element pe24_6(.reset(effective_rst), .clk(clk),  .in_a(a24_5to24_6), .in_b(b23_6to24_6),  .out_a(a24_6to24_7), .out_b(b24_6to25_6), .out_c(matrixC24_6));
processing_element pe24_7(.reset(effective_rst), .clk(clk),  .in_a(a24_6to24_7), .in_b(b23_7to24_7),  .out_a(a24_7to24_8), .out_b(b24_7to25_7), .out_c(matrixC24_7));
processing_element pe24_8(.reset(effective_rst), .clk(clk),  .in_a(a24_7to24_8), .in_b(b23_8to24_8),  .out_a(a24_8to24_9), .out_b(b24_8to25_8), .out_c(matrixC24_8));
processing_element pe24_9(.reset(effective_rst), .clk(clk),  .in_a(a24_8to24_9), .in_b(b23_9to24_9),  .out_a(a24_9to24_10), .out_b(b24_9to25_9), .out_c(matrixC24_9));
processing_element pe24_10(.reset(effective_rst), .clk(clk),  .in_a(a24_9to24_10), .in_b(b23_10to24_10),  .out_a(a24_10to24_11), .out_b(b24_10to25_10), .out_c(matrixC24_10));
processing_element pe24_11(.reset(effective_rst), .clk(clk),  .in_a(a24_10to24_11), .in_b(b23_11to24_11),  .out_a(a24_11to24_12), .out_b(b24_11to25_11), .out_c(matrixC24_11));
processing_element pe24_12(.reset(effective_rst), .clk(clk),  .in_a(a24_11to24_12), .in_b(b23_12to24_12),  .out_a(a24_12to24_13), .out_b(b24_12to25_12), .out_c(matrixC24_12));
processing_element pe24_13(.reset(effective_rst), .clk(clk),  .in_a(a24_12to24_13), .in_b(b23_13to24_13),  .out_a(a24_13to24_14), .out_b(b24_13to25_13), .out_c(matrixC24_13));
processing_element pe24_14(.reset(effective_rst), .clk(clk),  .in_a(a24_13to24_14), .in_b(b23_14to24_14),  .out_a(a24_14to24_15), .out_b(b24_14to25_14), .out_c(matrixC24_14));
processing_element pe24_15(.reset(effective_rst), .clk(clk),  .in_a(a24_14to24_15), .in_b(b23_15to24_15),  .out_a(a24_15to24_16), .out_b(b24_15to25_15), .out_c(matrixC24_15));
processing_element pe24_16(.reset(effective_rst), .clk(clk),  .in_a(a24_15to24_16), .in_b(b23_16to24_16),  .out_a(a24_16to24_17), .out_b(b24_16to25_16), .out_c(matrixC24_16));
processing_element pe24_17(.reset(effective_rst), .clk(clk),  .in_a(a24_16to24_17), .in_b(b23_17to24_17),  .out_a(a24_17to24_18), .out_b(b24_17to25_17), .out_c(matrixC24_17));
processing_element pe24_18(.reset(effective_rst), .clk(clk),  .in_a(a24_17to24_18), .in_b(b23_18to24_18),  .out_a(a24_18to24_19), .out_b(b24_18to25_18), .out_c(matrixC24_18));
processing_element pe24_19(.reset(effective_rst), .clk(clk),  .in_a(a24_18to24_19), .in_b(b23_19to24_19),  .out_a(a24_19to24_20), .out_b(b24_19to25_19), .out_c(matrixC24_19));
processing_element pe24_20(.reset(effective_rst), .clk(clk),  .in_a(a24_19to24_20), .in_b(b23_20to24_20),  .out_a(a24_20to24_21), .out_b(b24_20to25_20), .out_c(matrixC24_20));
processing_element pe24_21(.reset(effective_rst), .clk(clk),  .in_a(a24_20to24_21), .in_b(b23_21to24_21),  .out_a(a24_21to24_22), .out_b(b24_21to25_21), .out_c(matrixC24_21));
processing_element pe24_22(.reset(effective_rst), .clk(clk),  .in_a(a24_21to24_22), .in_b(b23_22to24_22),  .out_a(a24_22to24_23), .out_b(b24_22to25_22), .out_c(matrixC24_22));
processing_element pe24_23(.reset(effective_rst), .clk(clk),  .in_a(a24_22to24_23), .in_b(b23_23to24_23),  .out_a(a24_23to24_24), .out_b(b24_23to25_23), .out_c(matrixC24_23));
processing_element pe24_24(.reset(effective_rst), .clk(clk),  .in_a(a24_23to24_24), .in_b(b23_24to24_24),  .out_a(a24_24to24_25), .out_b(b24_24to25_24), .out_c(matrixC24_24));
processing_element pe24_25(.reset(effective_rst), .clk(clk),  .in_a(a24_24to24_25), .in_b(b23_25to24_25),  .out_a(a24_25to24_26), .out_b(b24_25to25_25), .out_c(matrixC24_25));
processing_element pe24_26(.reset(effective_rst), .clk(clk),  .in_a(a24_25to24_26), .in_b(b23_26to24_26),  .out_a(a24_26to24_27), .out_b(b24_26to25_26), .out_c(matrixC24_26));
processing_element pe24_27(.reset(effective_rst), .clk(clk),  .in_a(a24_26to24_27), .in_b(b23_27to24_27),  .out_a(a24_27to24_28), .out_b(b24_27to25_27), .out_c(matrixC24_27));
processing_element pe24_28(.reset(effective_rst), .clk(clk),  .in_a(a24_27to24_28), .in_b(b23_28to24_28),  .out_a(a24_28to24_29), .out_b(b24_28to25_28), .out_c(matrixC24_28));
processing_element pe24_29(.reset(effective_rst), .clk(clk),  .in_a(a24_28to24_29), .in_b(b23_29to24_29),  .out_a(a24_29to24_30), .out_b(b24_29to25_29), .out_c(matrixC24_29));
processing_element pe24_30(.reset(effective_rst), .clk(clk),  .in_a(a24_29to24_30), .in_b(b23_30to24_30),  .out_a(a24_30to24_31), .out_b(b24_30to25_30), .out_c(matrixC24_30));
processing_element pe24_31(.reset(effective_rst), .clk(clk),  .in_a(a24_30to24_31), .in_b(b23_31to24_31),  .out_a(a24_31to24_32), .out_b(b24_31to25_31), .out_c(matrixC24_31));
processing_element pe25_1(.reset(effective_rst), .clk(clk),  .in_a(a25_0to25_1), .in_b(b24_1to25_1),  .out_a(a25_1to25_2), .out_b(b25_1to26_1), .out_c(matrixC25_1));
processing_element pe25_2(.reset(effective_rst), .clk(clk),  .in_a(a25_1to25_2), .in_b(b24_2to25_2),  .out_a(a25_2to25_3), .out_b(b25_2to26_2), .out_c(matrixC25_2));
processing_element pe25_3(.reset(effective_rst), .clk(clk),  .in_a(a25_2to25_3), .in_b(b24_3to25_3),  .out_a(a25_3to25_4), .out_b(b25_3to26_3), .out_c(matrixC25_3));
processing_element pe25_4(.reset(effective_rst), .clk(clk),  .in_a(a25_3to25_4), .in_b(b24_4to25_4),  .out_a(a25_4to25_5), .out_b(b25_4to26_4), .out_c(matrixC25_4));
processing_element pe25_5(.reset(effective_rst), .clk(clk),  .in_a(a25_4to25_5), .in_b(b24_5to25_5),  .out_a(a25_5to25_6), .out_b(b25_5to26_5), .out_c(matrixC25_5));
processing_element pe25_6(.reset(effective_rst), .clk(clk),  .in_a(a25_5to25_6), .in_b(b24_6to25_6),  .out_a(a25_6to25_7), .out_b(b25_6to26_6), .out_c(matrixC25_6));
processing_element pe25_7(.reset(effective_rst), .clk(clk),  .in_a(a25_6to25_7), .in_b(b24_7to25_7),  .out_a(a25_7to25_8), .out_b(b25_7to26_7), .out_c(matrixC25_7));
processing_element pe25_8(.reset(effective_rst), .clk(clk),  .in_a(a25_7to25_8), .in_b(b24_8to25_8),  .out_a(a25_8to25_9), .out_b(b25_8to26_8), .out_c(matrixC25_8));
processing_element pe25_9(.reset(effective_rst), .clk(clk),  .in_a(a25_8to25_9), .in_b(b24_9to25_9),  .out_a(a25_9to25_10), .out_b(b25_9to26_9), .out_c(matrixC25_9));
processing_element pe25_10(.reset(effective_rst), .clk(clk),  .in_a(a25_9to25_10), .in_b(b24_10to25_10),  .out_a(a25_10to25_11), .out_b(b25_10to26_10), .out_c(matrixC25_10));
processing_element pe25_11(.reset(effective_rst), .clk(clk),  .in_a(a25_10to25_11), .in_b(b24_11to25_11),  .out_a(a25_11to25_12), .out_b(b25_11to26_11), .out_c(matrixC25_11));
processing_element pe25_12(.reset(effective_rst), .clk(clk),  .in_a(a25_11to25_12), .in_b(b24_12to25_12),  .out_a(a25_12to25_13), .out_b(b25_12to26_12), .out_c(matrixC25_12));
processing_element pe25_13(.reset(effective_rst), .clk(clk),  .in_a(a25_12to25_13), .in_b(b24_13to25_13),  .out_a(a25_13to25_14), .out_b(b25_13to26_13), .out_c(matrixC25_13));
processing_element pe25_14(.reset(effective_rst), .clk(clk),  .in_a(a25_13to25_14), .in_b(b24_14to25_14),  .out_a(a25_14to25_15), .out_b(b25_14to26_14), .out_c(matrixC25_14));
processing_element pe25_15(.reset(effective_rst), .clk(clk),  .in_a(a25_14to25_15), .in_b(b24_15to25_15),  .out_a(a25_15to25_16), .out_b(b25_15to26_15), .out_c(matrixC25_15));
processing_element pe25_16(.reset(effective_rst), .clk(clk),  .in_a(a25_15to25_16), .in_b(b24_16to25_16),  .out_a(a25_16to25_17), .out_b(b25_16to26_16), .out_c(matrixC25_16));
processing_element pe25_17(.reset(effective_rst), .clk(clk),  .in_a(a25_16to25_17), .in_b(b24_17to25_17),  .out_a(a25_17to25_18), .out_b(b25_17to26_17), .out_c(matrixC25_17));
processing_element pe25_18(.reset(effective_rst), .clk(clk),  .in_a(a25_17to25_18), .in_b(b24_18to25_18),  .out_a(a25_18to25_19), .out_b(b25_18to26_18), .out_c(matrixC25_18));
processing_element pe25_19(.reset(effective_rst), .clk(clk),  .in_a(a25_18to25_19), .in_b(b24_19to25_19),  .out_a(a25_19to25_20), .out_b(b25_19to26_19), .out_c(matrixC25_19));
processing_element pe25_20(.reset(effective_rst), .clk(clk),  .in_a(a25_19to25_20), .in_b(b24_20to25_20),  .out_a(a25_20to25_21), .out_b(b25_20to26_20), .out_c(matrixC25_20));
processing_element pe25_21(.reset(effective_rst), .clk(clk),  .in_a(a25_20to25_21), .in_b(b24_21to25_21),  .out_a(a25_21to25_22), .out_b(b25_21to26_21), .out_c(matrixC25_21));
processing_element pe25_22(.reset(effective_rst), .clk(clk),  .in_a(a25_21to25_22), .in_b(b24_22to25_22),  .out_a(a25_22to25_23), .out_b(b25_22to26_22), .out_c(matrixC25_22));
processing_element pe25_23(.reset(effective_rst), .clk(clk),  .in_a(a25_22to25_23), .in_b(b24_23to25_23),  .out_a(a25_23to25_24), .out_b(b25_23to26_23), .out_c(matrixC25_23));
processing_element pe25_24(.reset(effective_rst), .clk(clk),  .in_a(a25_23to25_24), .in_b(b24_24to25_24),  .out_a(a25_24to25_25), .out_b(b25_24to26_24), .out_c(matrixC25_24));
processing_element pe25_25(.reset(effective_rst), .clk(clk),  .in_a(a25_24to25_25), .in_b(b24_25to25_25),  .out_a(a25_25to25_26), .out_b(b25_25to26_25), .out_c(matrixC25_25));
processing_element pe25_26(.reset(effective_rst), .clk(clk),  .in_a(a25_25to25_26), .in_b(b24_26to25_26),  .out_a(a25_26to25_27), .out_b(b25_26to26_26), .out_c(matrixC25_26));
processing_element pe25_27(.reset(effective_rst), .clk(clk),  .in_a(a25_26to25_27), .in_b(b24_27to25_27),  .out_a(a25_27to25_28), .out_b(b25_27to26_27), .out_c(matrixC25_27));
processing_element pe25_28(.reset(effective_rst), .clk(clk),  .in_a(a25_27to25_28), .in_b(b24_28to25_28),  .out_a(a25_28to25_29), .out_b(b25_28to26_28), .out_c(matrixC25_28));
processing_element pe25_29(.reset(effective_rst), .clk(clk),  .in_a(a25_28to25_29), .in_b(b24_29to25_29),  .out_a(a25_29to25_30), .out_b(b25_29to26_29), .out_c(matrixC25_29));
processing_element pe25_30(.reset(effective_rst), .clk(clk),  .in_a(a25_29to25_30), .in_b(b24_30to25_30),  .out_a(a25_30to25_31), .out_b(b25_30to26_30), .out_c(matrixC25_30));
processing_element pe25_31(.reset(effective_rst), .clk(clk),  .in_a(a25_30to25_31), .in_b(b24_31to25_31),  .out_a(a25_31to25_32), .out_b(b25_31to26_31), .out_c(matrixC25_31));
processing_element pe26_1(.reset(effective_rst), .clk(clk),  .in_a(a26_0to26_1), .in_b(b25_1to26_1),  .out_a(a26_1to26_2), .out_b(b26_1to27_1), .out_c(matrixC26_1));
processing_element pe26_2(.reset(effective_rst), .clk(clk),  .in_a(a26_1to26_2), .in_b(b25_2to26_2),  .out_a(a26_2to26_3), .out_b(b26_2to27_2), .out_c(matrixC26_2));
processing_element pe26_3(.reset(effective_rst), .clk(clk),  .in_a(a26_2to26_3), .in_b(b25_3to26_3),  .out_a(a26_3to26_4), .out_b(b26_3to27_3), .out_c(matrixC26_3));
processing_element pe26_4(.reset(effective_rst), .clk(clk),  .in_a(a26_3to26_4), .in_b(b25_4to26_4),  .out_a(a26_4to26_5), .out_b(b26_4to27_4), .out_c(matrixC26_4));
processing_element pe26_5(.reset(effective_rst), .clk(clk),  .in_a(a26_4to26_5), .in_b(b25_5to26_5),  .out_a(a26_5to26_6), .out_b(b26_5to27_5), .out_c(matrixC26_5));
processing_element pe26_6(.reset(effective_rst), .clk(clk),  .in_a(a26_5to26_6), .in_b(b25_6to26_6),  .out_a(a26_6to26_7), .out_b(b26_6to27_6), .out_c(matrixC26_6));
processing_element pe26_7(.reset(effective_rst), .clk(clk),  .in_a(a26_6to26_7), .in_b(b25_7to26_7),  .out_a(a26_7to26_8), .out_b(b26_7to27_7), .out_c(matrixC26_7));
processing_element pe26_8(.reset(effective_rst), .clk(clk),  .in_a(a26_7to26_8), .in_b(b25_8to26_8),  .out_a(a26_8to26_9), .out_b(b26_8to27_8), .out_c(matrixC26_8));
processing_element pe26_9(.reset(effective_rst), .clk(clk),  .in_a(a26_8to26_9), .in_b(b25_9to26_9),  .out_a(a26_9to26_10), .out_b(b26_9to27_9), .out_c(matrixC26_9));
processing_element pe26_10(.reset(effective_rst), .clk(clk),  .in_a(a26_9to26_10), .in_b(b25_10to26_10),  .out_a(a26_10to26_11), .out_b(b26_10to27_10), .out_c(matrixC26_10));
processing_element pe26_11(.reset(effective_rst), .clk(clk),  .in_a(a26_10to26_11), .in_b(b25_11to26_11),  .out_a(a26_11to26_12), .out_b(b26_11to27_11), .out_c(matrixC26_11));
processing_element pe26_12(.reset(effective_rst), .clk(clk),  .in_a(a26_11to26_12), .in_b(b25_12to26_12),  .out_a(a26_12to26_13), .out_b(b26_12to27_12), .out_c(matrixC26_12));
processing_element pe26_13(.reset(effective_rst), .clk(clk),  .in_a(a26_12to26_13), .in_b(b25_13to26_13),  .out_a(a26_13to26_14), .out_b(b26_13to27_13), .out_c(matrixC26_13));
processing_element pe26_14(.reset(effective_rst), .clk(clk),  .in_a(a26_13to26_14), .in_b(b25_14to26_14),  .out_a(a26_14to26_15), .out_b(b26_14to27_14), .out_c(matrixC26_14));
processing_element pe26_15(.reset(effective_rst), .clk(clk),  .in_a(a26_14to26_15), .in_b(b25_15to26_15),  .out_a(a26_15to26_16), .out_b(b26_15to27_15), .out_c(matrixC26_15));
processing_element pe26_16(.reset(effective_rst), .clk(clk),  .in_a(a26_15to26_16), .in_b(b25_16to26_16),  .out_a(a26_16to26_17), .out_b(b26_16to27_16), .out_c(matrixC26_16));
processing_element pe26_17(.reset(effective_rst), .clk(clk),  .in_a(a26_16to26_17), .in_b(b25_17to26_17),  .out_a(a26_17to26_18), .out_b(b26_17to27_17), .out_c(matrixC26_17));
processing_element pe26_18(.reset(effective_rst), .clk(clk),  .in_a(a26_17to26_18), .in_b(b25_18to26_18),  .out_a(a26_18to26_19), .out_b(b26_18to27_18), .out_c(matrixC26_18));
processing_element pe26_19(.reset(effective_rst), .clk(clk),  .in_a(a26_18to26_19), .in_b(b25_19to26_19),  .out_a(a26_19to26_20), .out_b(b26_19to27_19), .out_c(matrixC26_19));
processing_element pe26_20(.reset(effective_rst), .clk(clk),  .in_a(a26_19to26_20), .in_b(b25_20to26_20),  .out_a(a26_20to26_21), .out_b(b26_20to27_20), .out_c(matrixC26_20));
processing_element pe26_21(.reset(effective_rst), .clk(clk),  .in_a(a26_20to26_21), .in_b(b25_21to26_21),  .out_a(a26_21to26_22), .out_b(b26_21to27_21), .out_c(matrixC26_21));
processing_element pe26_22(.reset(effective_rst), .clk(clk),  .in_a(a26_21to26_22), .in_b(b25_22to26_22),  .out_a(a26_22to26_23), .out_b(b26_22to27_22), .out_c(matrixC26_22));
processing_element pe26_23(.reset(effective_rst), .clk(clk),  .in_a(a26_22to26_23), .in_b(b25_23to26_23),  .out_a(a26_23to26_24), .out_b(b26_23to27_23), .out_c(matrixC26_23));
processing_element pe26_24(.reset(effective_rst), .clk(clk),  .in_a(a26_23to26_24), .in_b(b25_24to26_24),  .out_a(a26_24to26_25), .out_b(b26_24to27_24), .out_c(matrixC26_24));
processing_element pe26_25(.reset(effective_rst), .clk(clk),  .in_a(a26_24to26_25), .in_b(b25_25to26_25),  .out_a(a26_25to26_26), .out_b(b26_25to27_25), .out_c(matrixC26_25));
processing_element pe26_26(.reset(effective_rst), .clk(clk),  .in_a(a26_25to26_26), .in_b(b25_26to26_26),  .out_a(a26_26to26_27), .out_b(b26_26to27_26), .out_c(matrixC26_26));
processing_element pe26_27(.reset(effective_rst), .clk(clk),  .in_a(a26_26to26_27), .in_b(b25_27to26_27),  .out_a(a26_27to26_28), .out_b(b26_27to27_27), .out_c(matrixC26_27));
processing_element pe26_28(.reset(effective_rst), .clk(clk),  .in_a(a26_27to26_28), .in_b(b25_28to26_28),  .out_a(a26_28to26_29), .out_b(b26_28to27_28), .out_c(matrixC26_28));
processing_element pe26_29(.reset(effective_rst), .clk(clk),  .in_a(a26_28to26_29), .in_b(b25_29to26_29),  .out_a(a26_29to26_30), .out_b(b26_29to27_29), .out_c(matrixC26_29));
processing_element pe26_30(.reset(effective_rst), .clk(clk),  .in_a(a26_29to26_30), .in_b(b25_30to26_30),  .out_a(a26_30to26_31), .out_b(b26_30to27_30), .out_c(matrixC26_30));
processing_element pe26_31(.reset(effective_rst), .clk(clk),  .in_a(a26_30to26_31), .in_b(b25_31to26_31),  .out_a(a26_31to26_32), .out_b(b26_31to27_31), .out_c(matrixC26_31));
processing_element pe27_1(.reset(effective_rst), .clk(clk),  .in_a(a27_0to27_1), .in_b(b26_1to27_1),  .out_a(a27_1to27_2), .out_b(b27_1to28_1), .out_c(matrixC27_1));
processing_element pe27_2(.reset(effective_rst), .clk(clk),  .in_a(a27_1to27_2), .in_b(b26_2to27_2),  .out_a(a27_2to27_3), .out_b(b27_2to28_2), .out_c(matrixC27_2));
processing_element pe27_3(.reset(effective_rst), .clk(clk),  .in_a(a27_2to27_3), .in_b(b26_3to27_3),  .out_a(a27_3to27_4), .out_b(b27_3to28_3), .out_c(matrixC27_3));
processing_element pe27_4(.reset(effective_rst), .clk(clk),  .in_a(a27_3to27_4), .in_b(b26_4to27_4),  .out_a(a27_4to27_5), .out_b(b27_4to28_4), .out_c(matrixC27_4));
processing_element pe27_5(.reset(effective_rst), .clk(clk),  .in_a(a27_4to27_5), .in_b(b26_5to27_5),  .out_a(a27_5to27_6), .out_b(b27_5to28_5), .out_c(matrixC27_5));
processing_element pe27_6(.reset(effective_rst), .clk(clk),  .in_a(a27_5to27_6), .in_b(b26_6to27_6),  .out_a(a27_6to27_7), .out_b(b27_6to28_6), .out_c(matrixC27_6));
processing_element pe27_7(.reset(effective_rst), .clk(clk),  .in_a(a27_6to27_7), .in_b(b26_7to27_7),  .out_a(a27_7to27_8), .out_b(b27_7to28_7), .out_c(matrixC27_7));
processing_element pe27_8(.reset(effective_rst), .clk(clk),  .in_a(a27_7to27_8), .in_b(b26_8to27_8),  .out_a(a27_8to27_9), .out_b(b27_8to28_8), .out_c(matrixC27_8));
processing_element pe27_9(.reset(effective_rst), .clk(clk),  .in_a(a27_8to27_9), .in_b(b26_9to27_9),  .out_a(a27_9to27_10), .out_b(b27_9to28_9), .out_c(matrixC27_9));
processing_element pe27_10(.reset(effective_rst), .clk(clk),  .in_a(a27_9to27_10), .in_b(b26_10to27_10),  .out_a(a27_10to27_11), .out_b(b27_10to28_10), .out_c(matrixC27_10));
processing_element pe27_11(.reset(effective_rst), .clk(clk),  .in_a(a27_10to27_11), .in_b(b26_11to27_11),  .out_a(a27_11to27_12), .out_b(b27_11to28_11), .out_c(matrixC27_11));
processing_element pe27_12(.reset(effective_rst), .clk(clk),  .in_a(a27_11to27_12), .in_b(b26_12to27_12),  .out_a(a27_12to27_13), .out_b(b27_12to28_12), .out_c(matrixC27_12));
processing_element pe27_13(.reset(effective_rst), .clk(clk),  .in_a(a27_12to27_13), .in_b(b26_13to27_13),  .out_a(a27_13to27_14), .out_b(b27_13to28_13), .out_c(matrixC27_13));
processing_element pe27_14(.reset(effective_rst), .clk(clk),  .in_a(a27_13to27_14), .in_b(b26_14to27_14),  .out_a(a27_14to27_15), .out_b(b27_14to28_14), .out_c(matrixC27_14));
processing_element pe27_15(.reset(effective_rst), .clk(clk),  .in_a(a27_14to27_15), .in_b(b26_15to27_15),  .out_a(a27_15to27_16), .out_b(b27_15to28_15), .out_c(matrixC27_15));
processing_element pe27_16(.reset(effective_rst), .clk(clk),  .in_a(a27_15to27_16), .in_b(b26_16to27_16),  .out_a(a27_16to27_17), .out_b(b27_16to28_16), .out_c(matrixC27_16));
processing_element pe27_17(.reset(effective_rst), .clk(clk),  .in_a(a27_16to27_17), .in_b(b26_17to27_17),  .out_a(a27_17to27_18), .out_b(b27_17to28_17), .out_c(matrixC27_17));
processing_element pe27_18(.reset(effective_rst), .clk(clk),  .in_a(a27_17to27_18), .in_b(b26_18to27_18),  .out_a(a27_18to27_19), .out_b(b27_18to28_18), .out_c(matrixC27_18));
processing_element pe27_19(.reset(effective_rst), .clk(clk),  .in_a(a27_18to27_19), .in_b(b26_19to27_19),  .out_a(a27_19to27_20), .out_b(b27_19to28_19), .out_c(matrixC27_19));
processing_element pe27_20(.reset(effective_rst), .clk(clk),  .in_a(a27_19to27_20), .in_b(b26_20to27_20),  .out_a(a27_20to27_21), .out_b(b27_20to28_20), .out_c(matrixC27_20));
processing_element pe27_21(.reset(effective_rst), .clk(clk),  .in_a(a27_20to27_21), .in_b(b26_21to27_21),  .out_a(a27_21to27_22), .out_b(b27_21to28_21), .out_c(matrixC27_21));
processing_element pe27_22(.reset(effective_rst), .clk(clk),  .in_a(a27_21to27_22), .in_b(b26_22to27_22),  .out_a(a27_22to27_23), .out_b(b27_22to28_22), .out_c(matrixC27_22));
processing_element pe27_23(.reset(effective_rst), .clk(clk),  .in_a(a27_22to27_23), .in_b(b26_23to27_23),  .out_a(a27_23to27_24), .out_b(b27_23to28_23), .out_c(matrixC27_23));
processing_element pe27_24(.reset(effective_rst), .clk(clk),  .in_a(a27_23to27_24), .in_b(b26_24to27_24),  .out_a(a27_24to27_25), .out_b(b27_24to28_24), .out_c(matrixC27_24));
processing_element pe27_25(.reset(effective_rst), .clk(clk),  .in_a(a27_24to27_25), .in_b(b26_25to27_25),  .out_a(a27_25to27_26), .out_b(b27_25to28_25), .out_c(matrixC27_25));
processing_element pe27_26(.reset(effective_rst), .clk(clk),  .in_a(a27_25to27_26), .in_b(b26_26to27_26),  .out_a(a27_26to27_27), .out_b(b27_26to28_26), .out_c(matrixC27_26));
processing_element pe27_27(.reset(effective_rst), .clk(clk),  .in_a(a27_26to27_27), .in_b(b26_27to27_27),  .out_a(a27_27to27_28), .out_b(b27_27to28_27), .out_c(matrixC27_27));
processing_element pe27_28(.reset(effective_rst), .clk(clk),  .in_a(a27_27to27_28), .in_b(b26_28to27_28),  .out_a(a27_28to27_29), .out_b(b27_28to28_28), .out_c(matrixC27_28));
processing_element pe27_29(.reset(effective_rst), .clk(clk),  .in_a(a27_28to27_29), .in_b(b26_29to27_29),  .out_a(a27_29to27_30), .out_b(b27_29to28_29), .out_c(matrixC27_29));
processing_element pe27_30(.reset(effective_rst), .clk(clk),  .in_a(a27_29to27_30), .in_b(b26_30to27_30),  .out_a(a27_30to27_31), .out_b(b27_30to28_30), .out_c(matrixC27_30));
processing_element pe27_31(.reset(effective_rst), .clk(clk),  .in_a(a27_30to27_31), .in_b(b26_31to27_31),  .out_a(a27_31to27_32), .out_b(b27_31to28_31), .out_c(matrixC27_31));
processing_element pe28_1(.reset(effective_rst), .clk(clk),  .in_a(a28_0to28_1), .in_b(b27_1to28_1),  .out_a(a28_1to28_2), .out_b(b28_1to29_1), .out_c(matrixC28_1));
processing_element pe28_2(.reset(effective_rst), .clk(clk),  .in_a(a28_1to28_2), .in_b(b27_2to28_2),  .out_a(a28_2to28_3), .out_b(b28_2to29_2), .out_c(matrixC28_2));
processing_element pe28_3(.reset(effective_rst), .clk(clk),  .in_a(a28_2to28_3), .in_b(b27_3to28_3),  .out_a(a28_3to28_4), .out_b(b28_3to29_3), .out_c(matrixC28_3));
processing_element pe28_4(.reset(effective_rst), .clk(clk),  .in_a(a28_3to28_4), .in_b(b27_4to28_4),  .out_a(a28_4to28_5), .out_b(b28_4to29_4), .out_c(matrixC28_4));
processing_element pe28_5(.reset(effective_rst), .clk(clk),  .in_a(a28_4to28_5), .in_b(b27_5to28_5),  .out_a(a28_5to28_6), .out_b(b28_5to29_5), .out_c(matrixC28_5));
processing_element pe28_6(.reset(effective_rst), .clk(clk),  .in_a(a28_5to28_6), .in_b(b27_6to28_6),  .out_a(a28_6to28_7), .out_b(b28_6to29_6), .out_c(matrixC28_6));
processing_element pe28_7(.reset(effective_rst), .clk(clk),  .in_a(a28_6to28_7), .in_b(b27_7to28_7),  .out_a(a28_7to28_8), .out_b(b28_7to29_7), .out_c(matrixC28_7));
processing_element pe28_8(.reset(effective_rst), .clk(clk),  .in_a(a28_7to28_8), .in_b(b27_8to28_8),  .out_a(a28_8to28_9), .out_b(b28_8to29_8), .out_c(matrixC28_8));
processing_element pe28_9(.reset(effective_rst), .clk(clk),  .in_a(a28_8to28_9), .in_b(b27_9to28_9),  .out_a(a28_9to28_10), .out_b(b28_9to29_9), .out_c(matrixC28_9));
processing_element pe28_10(.reset(effective_rst), .clk(clk),  .in_a(a28_9to28_10), .in_b(b27_10to28_10),  .out_a(a28_10to28_11), .out_b(b28_10to29_10), .out_c(matrixC28_10));
processing_element pe28_11(.reset(effective_rst), .clk(clk),  .in_a(a28_10to28_11), .in_b(b27_11to28_11),  .out_a(a28_11to28_12), .out_b(b28_11to29_11), .out_c(matrixC28_11));
processing_element pe28_12(.reset(effective_rst), .clk(clk),  .in_a(a28_11to28_12), .in_b(b27_12to28_12),  .out_a(a28_12to28_13), .out_b(b28_12to29_12), .out_c(matrixC28_12));
processing_element pe28_13(.reset(effective_rst), .clk(clk),  .in_a(a28_12to28_13), .in_b(b27_13to28_13),  .out_a(a28_13to28_14), .out_b(b28_13to29_13), .out_c(matrixC28_13));
processing_element pe28_14(.reset(effective_rst), .clk(clk),  .in_a(a28_13to28_14), .in_b(b27_14to28_14),  .out_a(a28_14to28_15), .out_b(b28_14to29_14), .out_c(matrixC28_14));
processing_element pe28_15(.reset(effective_rst), .clk(clk),  .in_a(a28_14to28_15), .in_b(b27_15to28_15),  .out_a(a28_15to28_16), .out_b(b28_15to29_15), .out_c(matrixC28_15));
processing_element pe28_16(.reset(effective_rst), .clk(clk),  .in_a(a28_15to28_16), .in_b(b27_16to28_16),  .out_a(a28_16to28_17), .out_b(b28_16to29_16), .out_c(matrixC28_16));
processing_element pe28_17(.reset(effective_rst), .clk(clk),  .in_a(a28_16to28_17), .in_b(b27_17to28_17),  .out_a(a28_17to28_18), .out_b(b28_17to29_17), .out_c(matrixC28_17));
processing_element pe28_18(.reset(effective_rst), .clk(clk),  .in_a(a28_17to28_18), .in_b(b27_18to28_18),  .out_a(a28_18to28_19), .out_b(b28_18to29_18), .out_c(matrixC28_18));
processing_element pe28_19(.reset(effective_rst), .clk(clk),  .in_a(a28_18to28_19), .in_b(b27_19to28_19),  .out_a(a28_19to28_20), .out_b(b28_19to29_19), .out_c(matrixC28_19));
processing_element pe28_20(.reset(effective_rst), .clk(clk),  .in_a(a28_19to28_20), .in_b(b27_20to28_20),  .out_a(a28_20to28_21), .out_b(b28_20to29_20), .out_c(matrixC28_20));
processing_element pe28_21(.reset(effective_rst), .clk(clk),  .in_a(a28_20to28_21), .in_b(b27_21to28_21),  .out_a(a28_21to28_22), .out_b(b28_21to29_21), .out_c(matrixC28_21));
processing_element pe28_22(.reset(effective_rst), .clk(clk),  .in_a(a28_21to28_22), .in_b(b27_22to28_22),  .out_a(a28_22to28_23), .out_b(b28_22to29_22), .out_c(matrixC28_22));
processing_element pe28_23(.reset(effective_rst), .clk(clk),  .in_a(a28_22to28_23), .in_b(b27_23to28_23),  .out_a(a28_23to28_24), .out_b(b28_23to29_23), .out_c(matrixC28_23));
processing_element pe28_24(.reset(effective_rst), .clk(clk),  .in_a(a28_23to28_24), .in_b(b27_24to28_24),  .out_a(a28_24to28_25), .out_b(b28_24to29_24), .out_c(matrixC28_24));
processing_element pe28_25(.reset(effective_rst), .clk(clk),  .in_a(a28_24to28_25), .in_b(b27_25to28_25),  .out_a(a28_25to28_26), .out_b(b28_25to29_25), .out_c(matrixC28_25));
processing_element pe28_26(.reset(effective_rst), .clk(clk),  .in_a(a28_25to28_26), .in_b(b27_26to28_26),  .out_a(a28_26to28_27), .out_b(b28_26to29_26), .out_c(matrixC28_26));
processing_element pe28_27(.reset(effective_rst), .clk(clk),  .in_a(a28_26to28_27), .in_b(b27_27to28_27),  .out_a(a28_27to28_28), .out_b(b28_27to29_27), .out_c(matrixC28_27));
processing_element pe28_28(.reset(effective_rst), .clk(clk),  .in_a(a28_27to28_28), .in_b(b27_28to28_28),  .out_a(a28_28to28_29), .out_b(b28_28to29_28), .out_c(matrixC28_28));
processing_element pe28_29(.reset(effective_rst), .clk(clk),  .in_a(a28_28to28_29), .in_b(b27_29to28_29),  .out_a(a28_29to28_30), .out_b(b28_29to29_29), .out_c(matrixC28_29));
processing_element pe28_30(.reset(effective_rst), .clk(clk),  .in_a(a28_29to28_30), .in_b(b27_30to28_30),  .out_a(a28_30to28_31), .out_b(b28_30to29_30), .out_c(matrixC28_30));
processing_element pe28_31(.reset(effective_rst), .clk(clk),  .in_a(a28_30to28_31), .in_b(b27_31to28_31),  .out_a(a28_31to28_32), .out_b(b28_31to29_31), .out_c(matrixC28_31));
processing_element pe29_1(.reset(effective_rst), .clk(clk),  .in_a(a29_0to29_1), .in_b(b28_1to29_1),  .out_a(a29_1to29_2), .out_b(b29_1to30_1), .out_c(matrixC29_1));
processing_element pe29_2(.reset(effective_rst), .clk(clk),  .in_a(a29_1to29_2), .in_b(b28_2to29_2),  .out_a(a29_2to29_3), .out_b(b29_2to30_2), .out_c(matrixC29_2));
processing_element pe29_3(.reset(effective_rst), .clk(clk),  .in_a(a29_2to29_3), .in_b(b28_3to29_3),  .out_a(a29_3to29_4), .out_b(b29_3to30_3), .out_c(matrixC29_3));
processing_element pe29_4(.reset(effective_rst), .clk(clk),  .in_a(a29_3to29_4), .in_b(b28_4to29_4),  .out_a(a29_4to29_5), .out_b(b29_4to30_4), .out_c(matrixC29_4));
processing_element pe29_5(.reset(effective_rst), .clk(clk),  .in_a(a29_4to29_5), .in_b(b28_5to29_5),  .out_a(a29_5to29_6), .out_b(b29_5to30_5), .out_c(matrixC29_5));
processing_element pe29_6(.reset(effective_rst), .clk(clk),  .in_a(a29_5to29_6), .in_b(b28_6to29_6),  .out_a(a29_6to29_7), .out_b(b29_6to30_6), .out_c(matrixC29_6));
processing_element pe29_7(.reset(effective_rst), .clk(clk),  .in_a(a29_6to29_7), .in_b(b28_7to29_7),  .out_a(a29_7to29_8), .out_b(b29_7to30_7), .out_c(matrixC29_7));
processing_element pe29_8(.reset(effective_rst), .clk(clk),  .in_a(a29_7to29_8), .in_b(b28_8to29_8),  .out_a(a29_8to29_9), .out_b(b29_8to30_8), .out_c(matrixC29_8));
processing_element pe29_9(.reset(effective_rst), .clk(clk),  .in_a(a29_8to29_9), .in_b(b28_9to29_9),  .out_a(a29_9to29_10), .out_b(b29_9to30_9), .out_c(matrixC29_9));
processing_element pe29_10(.reset(effective_rst), .clk(clk),  .in_a(a29_9to29_10), .in_b(b28_10to29_10),  .out_a(a29_10to29_11), .out_b(b29_10to30_10), .out_c(matrixC29_10));
processing_element pe29_11(.reset(effective_rst), .clk(clk),  .in_a(a29_10to29_11), .in_b(b28_11to29_11),  .out_a(a29_11to29_12), .out_b(b29_11to30_11), .out_c(matrixC29_11));
processing_element pe29_12(.reset(effective_rst), .clk(clk),  .in_a(a29_11to29_12), .in_b(b28_12to29_12),  .out_a(a29_12to29_13), .out_b(b29_12to30_12), .out_c(matrixC29_12));
processing_element pe29_13(.reset(effective_rst), .clk(clk),  .in_a(a29_12to29_13), .in_b(b28_13to29_13),  .out_a(a29_13to29_14), .out_b(b29_13to30_13), .out_c(matrixC29_13));
processing_element pe29_14(.reset(effective_rst), .clk(clk),  .in_a(a29_13to29_14), .in_b(b28_14to29_14),  .out_a(a29_14to29_15), .out_b(b29_14to30_14), .out_c(matrixC29_14));
processing_element pe29_15(.reset(effective_rst), .clk(clk),  .in_a(a29_14to29_15), .in_b(b28_15to29_15),  .out_a(a29_15to29_16), .out_b(b29_15to30_15), .out_c(matrixC29_15));
processing_element pe29_16(.reset(effective_rst), .clk(clk),  .in_a(a29_15to29_16), .in_b(b28_16to29_16),  .out_a(a29_16to29_17), .out_b(b29_16to30_16), .out_c(matrixC29_16));
processing_element pe29_17(.reset(effective_rst), .clk(clk),  .in_a(a29_16to29_17), .in_b(b28_17to29_17),  .out_a(a29_17to29_18), .out_b(b29_17to30_17), .out_c(matrixC29_17));
processing_element pe29_18(.reset(effective_rst), .clk(clk),  .in_a(a29_17to29_18), .in_b(b28_18to29_18),  .out_a(a29_18to29_19), .out_b(b29_18to30_18), .out_c(matrixC29_18));
processing_element pe29_19(.reset(effective_rst), .clk(clk),  .in_a(a29_18to29_19), .in_b(b28_19to29_19),  .out_a(a29_19to29_20), .out_b(b29_19to30_19), .out_c(matrixC29_19));
processing_element pe29_20(.reset(effective_rst), .clk(clk),  .in_a(a29_19to29_20), .in_b(b28_20to29_20),  .out_a(a29_20to29_21), .out_b(b29_20to30_20), .out_c(matrixC29_20));
processing_element pe29_21(.reset(effective_rst), .clk(clk),  .in_a(a29_20to29_21), .in_b(b28_21to29_21),  .out_a(a29_21to29_22), .out_b(b29_21to30_21), .out_c(matrixC29_21));
processing_element pe29_22(.reset(effective_rst), .clk(clk),  .in_a(a29_21to29_22), .in_b(b28_22to29_22),  .out_a(a29_22to29_23), .out_b(b29_22to30_22), .out_c(matrixC29_22));
processing_element pe29_23(.reset(effective_rst), .clk(clk),  .in_a(a29_22to29_23), .in_b(b28_23to29_23),  .out_a(a29_23to29_24), .out_b(b29_23to30_23), .out_c(matrixC29_23));
processing_element pe29_24(.reset(effective_rst), .clk(clk),  .in_a(a29_23to29_24), .in_b(b28_24to29_24),  .out_a(a29_24to29_25), .out_b(b29_24to30_24), .out_c(matrixC29_24));
processing_element pe29_25(.reset(effective_rst), .clk(clk),  .in_a(a29_24to29_25), .in_b(b28_25to29_25),  .out_a(a29_25to29_26), .out_b(b29_25to30_25), .out_c(matrixC29_25));
processing_element pe29_26(.reset(effective_rst), .clk(clk),  .in_a(a29_25to29_26), .in_b(b28_26to29_26),  .out_a(a29_26to29_27), .out_b(b29_26to30_26), .out_c(matrixC29_26));
processing_element pe29_27(.reset(effective_rst), .clk(clk),  .in_a(a29_26to29_27), .in_b(b28_27to29_27),  .out_a(a29_27to29_28), .out_b(b29_27to30_27), .out_c(matrixC29_27));
processing_element pe29_28(.reset(effective_rst), .clk(clk),  .in_a(a29_27to29_28), .in_b(b28_28to29_28),  .out_a(a29_28to29_29), .out_b(b29_28to30_28), .out_c(matrixC29_28));
processing_element pe29_29(.reset(effective_rst), .clk(clk),  .in_a(a29_28to29_29), .in_b(b28_29to29_29),  .out_a(a29_29to29_30), .out_b(b29_29to30_29), .out_c(matrixC29_29));
processing_element pe29_30(.reset(effective_rst), .clk(clk),  .in_a(a29_29to29_30), .in_b(b28_30to29_30),  .out_a(a29_30to29_31), .out_b(b29_30to30_30), .out_c(matrixC29_30));
processing_element pe29_31(.reset(effective_rst), .clk(clk),  .in_a(a29_30to29_31), .in_b(b28_31to29_31),  .out_a(a29_31to29_32), .out_b(b29_31to30_31), .out_c(matrixC29_31));
processing_element pe30_1(.reset(effective_rst), .clk(clk),  .in_a(a30_0to30_1), .in_b(b29_1to30_1),  .out_a(a30_1to30_2), .out_b(b30_1to31_1), .out_c(matrixC30_1));
processing_element pe30_2(.reset(effective_rst), .clk(clk),  .in_a(a30_1to30_2), .in_b(b29_2to30_2),  .out_a(a30_2to30_3), .out_b(b30_2to31_2), .out_c(matrixC30_2));
processing_element pe30_3(.reset(effective_rst), .clk(clk),  .in_a(a30_2to30_3), .in_b(b29_3to30_3),  .out_a(a30_3to30_4), .out_b(b30_3to31_3), .out_c(matrixC30_3));
processing_element pe30_4(.reset(effective_rst), .clk(clk),  .in_a(a30_3to30_4), .in_b(b29_4to30_4),  .out_a(a30_4to30_5), .out_b(b30_4to31_4), .out_c(matrixC30_4));
processing_element pe30_5(.reset(effective_rst), .clk(clk),  .in_a(a30_4to30_5), .in_b(b29_5to30_5),  .out_a(a30_5to30_6), .out_b(b30_5to31_5), .out_c(matrixC30_5));
processing_element pe30_6(.reset(effective_rst), .clk(clk),  .in_a(a30_5to30_6), .in_b(b29_6to30_6),  .out_a(a30_6to30_7), .out_b(b30_6to31_6), .out_c(matrixC30_6));
processing_element pe30_7(.reset(effective_rst), .clk(clk),  .in_a(a30_6to30_7), .in_b(b29_7to30_7),  .out_a(a30_7to30_8), .out_b(b30_7to31_7), .out_c(matrixC30_7));
processing_element pe30_8(.reset(effective_rst), .clk(clk),  .in_a(a30_7to30_8), .in_b(b29_8to30_8),  .out_a(a30_8to30_9), .out_b(b30_8to31_8), .out_c(matrixC30_8));
processing_element pe30_9(.reset(effective_rst), .clk(clk),  .in_a(a30_8to30_9), .in_b(b29_9to30_9),  .out_a(a30_9to30_10), .out_b(b30_9to31_9), .out_c(matrixC30_9));
processing_element pe30_10(.reset(effective_rst), .clk(clk),  .in_a(a30_9to30_10), .in_b(b29_10to30_10),  .out_a(a30_10to30_11), .out_b(b30_10to31_10), .out_c(matrixC30_10));
processing_element pe30_11(.reset(effective_rst), .clk(clk),  .in_a(a30_10to30_11), .in_b(b29_11to30_11),  .out_a(a30_11to30_12), .out_b(b30_11to31_11), .out_c(matrixC30_11));
processing_element pe30_12(.reset(effective_rst), .clk(clk),  .in_a(a30_11to30_12), .in_b(b29_12to30_12),  .out_a(a30_12to30_13), .out_b(b30_12to31_12), .out_c(matrixC30_12));
processing_element pe30_13(.reset(effective_rst), .clk(clk),  .in_a(a30_12to30_13), .in_b(b29_13to30_13),  .out_a(a30_13to30_14), .out_b(b30_13to31_13), .out_c(matrixC30_13));
processing_element pe30_14(.reset(effective_rst), .clk(clk),  .in_a(a30_13to30_14), .in_b(b29_14to30_14),  .out_a(a30_14to30_15), .out_b(b30_14to31_14), .out_c(matrixC30_14));
processing_element pe30_15(.reset(effective_rst), .clk(clk),  .in_a(a30_14to30_15), .in_b(b29_15to30_15),  .out_a(a30_15to30_16), .out_b(b30_15to31_15), .out_c(matrixC30_15));
processing_element pe30_16(.reset(effective_rst), .clk(clk),  .in_a(a30_15to30_16), .in_b(b29_16to30_16),  .out_a(a30_16to30_17), .out_b(b30_16to31_16), .out_c(matrixC30_16));
processing_element pe30_17(.reset(effective_rst), .clk(clk),  .in_a(a30_16to30_17), .in_b(b29_17to30_17),  .out_a(a30_17to30_18), .out_b(b30_17to31_17), .out_c(matrixC30_17));
processing_element pe30_18(.reset(effective_rst), .clk(clk),  .in_a(a30_17to30_18), .in_b(b29_18to30_18),  .out_a(a30_18to30_19), .out_b(b30_18to31_18), .out_c(matrixC30_18));
processing_element pe30_19(.reset(effective_rst), .clk(clk),  .in_a(a30_18to30_19), .in_b(b29_19to30_19),  .out_a(a30_19to30_20), .out_b(b30_19to31_19), .out_c(matrixC30_19));
processing_element pe30_20(.reset(effective_rst), .clk(clk),  .in_a(a30_19to30_20), .in_b(b29_20to30_20),  .out_a(a30_20to30_21), .out_b(b30_20to31_20), .out_c(matrixC30_20));
processing_element pe30_21(.reset(effective_rst), .clk(clk),  .in_a(a30_20to30_21), .in_b(b29_21to30_21),  .out_a(a30_21to30_22), .out_b(b30_21to31_21), .out_c(matrixC30_21));
processing_element pe30_22(.reset(effective_rst), .clk(clk),  .in_a(a30_21to30_22), .in_b(b29_22to30_22),  .out_a(a30_22to30_23), .out_b(b30_22to31_22), .out_c(matrixC30_22));
processing_element pe30_23(.reset(effective_rst), .clk(clk),  .in_a(a30_22to30_23), .in_b(b29_23to30_23),  .out_a(a30_23to30_24), .out_b(b30_23to31_23), .out_c(matrixC30_23));
processing_element pe30_24(.reset(effective_rst), .clk(clk),  .in_a(a30_23to30_24), .in_b(b29_24to30_24),  .out_a(a30_24to30_25), .out_b(b30_24to31_24), .out_c(matrixC30_24));
processing_element pe30_25(.reset(effective_rst), .clk(clk),  .in_a(a30_24to30_25), .in_b(b29_25to30_25),  .out_a(a30_25to30_26), .out_b(b30_25to31_25), .out_c(matrixC30_25));
processing_element pe30_26(.reset(effective_rst), .clk(clk),  .in_a(a30_25to30_26), .in_b(b29_26to30_26),  .out_a(a30_26to30_27), .out_b(b30_26to31_26), .out_c(matrixC30_26));
processing_element pe30_27(.reset(effective_rst), .clk(clk),  .in_a(a30_26to30_27), .in_b(b29_27to30_27),  .out_a(a30_27to30_28), .out_b(b30_27to31_27), .out_c(matrixC30_27));
processing_element pe30_28(.reset(effective_rst), .clk(clk),  .in_a(a30_27to30_28), .in_b(b29_28to30_28),  .out_a(a30_28to30_29), .out_b(b30_28to31_28), .out_c(matrixC30_28));
processing_element pe30_29(.reset(effective_rst), .clk(clk),  .in_a(a30_28to30_29), .in_b(b29_29to30_29),  .out_a(a30_29to30_30), .out_b(b30_29to31_29), .out_c(matrixC30_29));
processing_element pe30_30(.reset(effective_rst), .clk(clk),  .in_a(a30_29to30_30), .in_b(b29_30to30_30),  .out_a(a30_30to30_31), .out_b(b30_30to31_30), .out_c(matrixC30_30));
processing_element pe30_31(.reset(effective_rst), .clk(clk),  .in_a(a30_30to30_31), .in_b(b29_31to30_31),  .out_a(a30_31to30_32), .out_b(b30_31to31_31), .out_c(matrixC30_31));
processing_element pe31_1(.reset(effective_rst), .clk(clk),  .in_a(a31_0to31_1), .in_b(b30_1to31_1),  .out_a(a31_1to31_2), .out_b(b31_1to32_1), .out_c(matrixC31_1));
processing_element pe31_2(.reset(effective_rst), .clk(clk),  .in_a(a31_1to31_2), .in_b(b30_2to31_2),  .out_a(a31_2to31_3), .out_b(b31_2to32_2), .out_c(matrixC31_2));
processing_element pe31_3(.reset(effective_rst), .clk(clk),  .in_a(a31_2to31_3), .in_b(b30_3to31_3),  .out_a(a31_3to31_4), .out_b(b31_3to32_3), .out_c(matrixC31_3));
processing_element pe31_4(.reset(effective_rst), .clk(clk),  .in_a(a31_3to31_4), .in_b(b30_4to31_4),  .out_a(a31_4to31_5), .out_b(b31_4to32_4), .out_c(matrixC31_4));
processing_element pe31_5(.reset(effective_rst), .clk(clk),  .in_a(a31_4to31_5), .in_b(b30_5to31_5),  .out_a(a31_5to31_6), .out_b(b31_5to32_5), .out_c(matrixC31_5));
processing_element pe31_6(.reset(effective_rst), .clk(clk),  .in_a(a31_5to31_6), .in_b(b30_6to31_6),  .out_a(a31_6to31_7), .out_b(b31_6to32_6), .out_c(matrixC31_6));
processing_element pe31_7(.reset(effective_rst), .clk(clk),  .in_a(a31_6to31_7), .in_b(b30_7to31_7),  .out_a(a31_7to31_8), .out_b(b31_7to32_7), .out_c(matrixC31_7));
processing_element pe31_8(.reset(effective_rst), .clk(clk),  .in_a(a31_7to31_8), .in_b(b30_8to31_8),  .out_a(a31_8to31_9), .out_b(b31_8to32_8), .out_c(matrixC31_8));
processing_element pe31_9(.reset(effective_rst), .clk(clk),  .in_a(a31_8to31_9), .in_b(b30_9to31_9),  .out_a(a31_9to31_10), .out_b(b31_9to32_9), .out_c(matrixC31_9));
processing_element pe31_10(.reset(effective_rst), .clk(clk),  .in_a(a31_9to31_10), .in_b(b30_10to31_10),  .out_a(a31_10to31_11), .out_b(b31_10to32_10), .out_c(matrixC31_10));
processing_element pe31_11(.reset(effective_rst), .clk(clk),  .in_a(a31_10to31_11), .in_b(b30_11to31_11),  .out_a(a31_11to31_12), .out_b(b31_11to32_11), .out_c(matrixC31_11));
processing_element pe31_12(.reset(effective_rst), .clk(clk),  .in_a(a31_11to31_12), .in_b(b30_12to31_12),  .out_a(a31_12to31_13), .out_b(b31_12to32_12), .out_c(matrixC31_12));
processing_element pe31_13(.reset(effective_rst), .clk(clk),  .in_a(a31_12to31_13), .in_b(b30_13to31_13),  .out_a(a31_13to31_14), .out_b(b31_13to32_13), .out_c(matrixC31_13));
processing_element pe31_14(.reset(effective_rst), .clk(clk),  .in_a(a31_13to31_14), .in_b(b30_14to31_14),  .out_a(a31_14to31_15), .out_b(b31_14to32_14), .out_c(matrixC31_14));
processing_element pe31_15(.reset(effective_rst), .clk(clk),  .in_a(a31_14to31_15), .in_b(b30_15to31_15),  .out_a(a31_15to31_16), .out_b(b31_15to32_15), .out_c(matrixC31_15));
processing_element pe31_16(.reset(effective_rst), .clk(clk),  .in_a(a31_15to31_16), .in_b(b30_16to31_16),  .out_a(a31_16to31_17), .out_b(b31_16to32_16), .out_c(matrixC31_16));
processing_element pe31_17(.reset(effective_rst), .clk(clk),  .in_a(a31_16to31_17), .in_b(b30_17to31_17),  .out_a(a31_17to31_18), .out_b(b31_17to32_17), .out_c(matrixC31_17));
processing_element pe31_18(.reset(effective_rst), .clk(clk),  .in_a(a31_17to31_18), .in_b(b30_18to31_18),  .out_a(a31_18to31_19), .out_b(b31_18to32_18), .out_c(matrixC31_18));
processing_element pe31_19(.reset(effective_rst), .clk(clk),  .in_a(a31_18to31_19), .in_b(b30_19to31_19),  .out_a(a31_19to31_20), .out_b(b31_19to32_19), .out_c(matrixC31_19));
processing_element pe31_20(.reset(effective_rst), .clk(clk),  .in_a(a31_19to31_20), .in_b(b30_20to31_20),  .out_a(a31_20to31_21), .out_b(b31_20to32_20), .out_c(matrixC31_20));
processing_element pe31_21(.reset(effective_rst), .clk(clk),  .in_a(a31_20to31_21), .in_b(b30_21to31_21),  .out_a(a31_21to31_22), .out_b(b31_21to32_21), .out_c(matrixC31_21));
processing_element pe31_22(.reset(effective_rst), .clk(clk),  .in_a(a31_21to31_22), .in_b(b30_22to31_22),  .out_a(a31_22to31_23), .out_b(b31_22to32_22), .out_c(matrixC31_22));
processing_element pe31_23(.reset(effective_rst), .clk(clk),  .in_a(a31_22to31_23), .in_b(b30_23to31_23),  .out_a(a31_23to31_24), .out_b(b31_23to32_23), .out_c(matrixC31_23));
processing_element pe31_24(.reset(effective_rst), .clk(clk),  .in_a(a31_23to31_24), .in_b(b30_24to31_24),  .out_a(a31_24to31_25), .out_b(b31_24to32_24), .out_c(matrixC31_24));
processing_element pe31_25(.reset(effective_rst), .clk(clk),  .in_a(a31_24to31_25), .in_b(b30_25to31_25),  .out_a(a31_25to31_26), .out_b(b31_25to32_25), .out_c(matrixC31_25));
processing_element pe31_26(.reset(effective_rst), .clk(clk),  .in_a(a31_25to31_26), .in_b(b30_26to31_26),  .out_a(a31_26to31_27), .out_b(b31_26to32_26), .out_c(matrixC31_26));
processing_element pe31_27(.reset(effective_rst), .clk(clk),  .in_a(a31_26to31_27), .in_b(b30_27to31_27),  .out_a(a31_27to31_28), .out_b(b31_27to32_27), .out_c(matrixC31_27));
processing_element pe31_28(.reset(effective_rst), .clk(clk),  .in_a(a31_27to31_28), .in_b(b30_28to31_28),  .out_a(a31_28to31_29), .out_b(b31_28to32_28), .out_c(matrixC31_28));
processing_element pe31_29(.reset(effective_rst), .clk(clk),  .in_a(a31_28to31_29), .in_b(b30_29to31_29),  .out_a(a31_29to31_30), .out_b(b31_29to32_29), .out_c(matrixC31_29));
processing_element pe31_30(.reset(effective_rst), .clk(clk),  .in_a(a31_29to31_30), .in_b(b30_30to31_30),  .out_a(a31_30to31_31), .out_b(b31_30to32_30), .out_c(matrixC31_30));
processing_element pe31_31(.reset(effective_rst), .clk(clk),  .in_a(a31_30to31_31), .in_b(b30_31to31_31),  .out_a(a31_31to31_32), .out_b(b31_31to32_31), .out_c(matrixC31_31));
assign a_data_out = {a31_31to31_32,a30_31to30_32,a29_31to29_32,a28_31to28_32,a27_31to27_32,a26_31to26_32,a25_31to25_32,a24_31to24_32,a23_31to23_32,a22_31to22_32,a21_31to21_32,a20_31to20_32,a19_31to19_32,a18_31to18_32,a17_31to17_32,a16_31to16_32,a15_31to15_32,a14_31to14_32,a13_31to13_32,a12_31to12_32,a11_31to11_32,a10_31to10_32,a9_31to9_32,a8_31to8_32,a7_31to7_32,a6_31to6_32,a5_31to5_32,a4_31to4_32,a3_31to3_32,a2_31to2_32,a1_31to1_32,a0_31to0_32};
assign b_data_out = {b31_31to32_31,b31_30to32_30,b31_29to32_29,b31_28to32_28,b31_27to32_27,b31_26to32_26,b31_25to32_25,b31_24to32_24,b31_23to32_23,b31_22to32_22,b31_21to32_21,b31_20to32_20,b31_19to32_19,b31_18to32_18,b31_17to32_17,b31_16to32_16,b31_15to32_15,b31_14to32_14,b31_13to32_13,b31_12to32_12,b31_11to32_11,b31_10to32_10,b31_9to32_9,b31_8to32_8,b31_7to32_7,b31_6to32_6,b31_5to32_5,b31_4to32_4,b31_3to32_3,b31_2to32_2,b31_1to32_1,b31_0to32_0};

endmodule

module processing_element(
 reset, 
 clk, 
 in_a,
 in_b, 
 out_a, 
 out_b, 
 out_c
 );

 input reset;
 input clk;
 input  [`DWIDTH-1:0] in_a;
 input  [`DWIDTH-1:0] in_b;
 output [`DWIDTH-1:0] out_a;
 output [`DWIDTH-1:0] out_b;
 output [`DWIDTH-1:0] out_c;  //reduced precision

 reg [`DWIDTH-1:0] out_a;
 reg [`DWIDTH-1:0] out_b;
 wire [`DWIDTH-1:0] out_c;

 wire [`DWIDTH-1:0] out_mac;

 assign out_c = out_mac;

 seq_mac u_mac(.a(in_a), .b(in_b), .out(out_mac), .reset(reset), .clk(clk));

 always @(posedge clk)begin
    if(reset) begin
      out_a<=0;
      out_b<=0;
    end
    else begin  
      out_a<=in_a;
      out_b<=in_b;
    end
 end
 
endmodule

module seq_mac(a, b, out, reset, clk);
input [`DWIDTH-1:0] a;
input [`DWIDTH-1:0] b;
input reset;
input clk;
output [`DWIDTH-1:0] out;

reg [`DWIDTH-1:0] out;
wire [`DWIDTH-1:0] mul_out;
wire [`DWIDTH-1:0] add_out;

reg [`DWIDTH-1:0] a_flopped;
reg [`DWIDTH-1:0] b_flopped;

wire [2*`DWIDTH-1:0] mul_out_temp;
reg [2*`DWIDTH-1:0] mul_out_temp_reg;

always @(posedge clk) begin
  if (reset) begin
    a_flopped <= 0;
    b_flopped <= 0;
  end else begin
    a_flopped <= a;
    b_flopped <= b;
  end
end

//assign mul_out = a * b;
qmult mult_u1(.i_multiplicand(a_flopped), .i_multiplier(b_flopped), .o_result(mul_out_temp));

always @(posedge clk) begin
  if (reset) begin
    mul_out_temp_reg <= 0;
  end else begin
    mul_out_temp_reg <= mul_out_temp;
  end
end

//down cast the result
assign mul_out = 
    (mul_out_temp_reg[2*`DWIDTH-1] == 0) ?  //positive number
        (
           (|(mul_out_temp_reg[2*`DWIDTH-2 : `DWIDTH-1])) ?  //is any bit from 14:7 is 1, that means overlfow
             {mul_out_temp_reg[2*`DWIDTH-1] , {(`DWIDTH-1){1'b1}}} : //sign bit and then all 1s
             {mul_out_temp_reg[2*`DWIDTH-1] , mul_out_temp_reg[`DWIDTH-2:0]} 
        )
        : //negative number
        (
           (|(mul_out_temp_reg[2*`DWIDTH-2 : `DWIDTH-1])) ?  //is any bit from 14:7 is 0, that means overlfow
             {mul_out_temp_reg[2*`DWIDTH-1] , mul_out_temp_reg[`DWIDTH-2:0]} :
             {mul_out_temp_reg[2*`DWIDTH-1] , {(`DWIDTH-1){1'b0}}} //sign bit and then all 0s
        );


//we just truncate the higher bits of the product
//assign add_out = mul_out + out;
qadd add_u1(.a(out), .b(mul_out), .c(add_out));

always @(posedge clk) begin
  if (reset) begin
    out <= 0;
  end else begin
    out <= add_out;
  end
end

endmodule

module qmult(i_multiplicand,i_multiplier,o_result);
input [`DWIDTH-1:0] i_multiplicand;
input [`DWIDTH-1:0] i_multiplier;
output [2*`DWIDTH-1:0] o_result;

assign o_result = i_multiplicand * i_multiplier;
//DW02_mult #(`DWIDTH,`DWIDTH) u_mult(.A(i_multiplicand), .B(i_multiplier), .TC(1'b1), .PRODUCT(o_result));

endmodule

module qadd(a,b,c);
input [`DWIDTH-1:0] a;
input [`DWIDTH-1:0] b;
output [`DWIDTH-1:0] c;

assign c = a + b;
//DW01_add #(`DWIDTH) u_add(.A(a), .B(b), .CI(1'b0), .SUM(c), .CO());
endmodule
