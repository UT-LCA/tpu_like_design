module conv_test();

task run();
begin
  initialize_brams();
  convolution_test();
  //compare_outputs();
end
endtask

integer a_start_addr = 0;
integer b_start_addr = 0;
integer c_start_addr = 200;

integer batch_size = 2;
integer inp_channels = 4;
integer out_channels = 4;
integer inp_height = 8;
integer inp_width = 8;
integer filter_height = 2;
integer filter_width = 2;

////////////////////////////////////////////
// Note: Data layout is NCHW
// This means that the fastest changing dimension
// is W. That is, as address increases, we first change
// W, then H, then C and then N.
////////////////////////////////////////////

////////////////////////////////////////////
// 4D input matrix
////////////////////////////////////////////

/*
>>> a = np.random.randint(low=0, high=3,size=(2,4,8,8), dtype=np.uint8)
>>> a
array([[[[1, 1, 1, 1, 1, 1, 2, 0],
         [0, 1, 1, 1, 1, 2, 2, 1],
         [0, 0, 0, 2, 2, 0, 0, 2],
         [1, 0, 0, 2, 2, 2, 0, 1],
         [2, 2, 2, 2, 0, 2, 1, 1],
         [2, 1, 1, 2, 2, 1, 0, 0],
         [0, 0, 0, 0, 0, 1, 2, 2],
         [0, 2, 0, 2, 1, 0, 2, 1]],

        [[0, 0, 0, 0, 0, 0, 1, 0],
         [1, 2, 1, 0, 1, 2, 1, 0],
         [1, 1, 2, 0, 0, 1, 0, 0],
         [2, 2, 2, 0, 2, 2, 1, 2],
         [1, 2, 0, 2, 1, 2, 1, 0],
         [2, 2, 0, 0, 0, 0, 1, 2],
         [1, 0, 2, 1, 1, 0, 1, 0],
         [1, 1, 0, 2, 0, 2, 1, 2]],

        [[0, 1, 2, 2, 1, 0, 2, 0],
         [2, 0, 1, 1, 2, 0, 0, 2],
         [1, 1, 1, 0, 1, 0, 1, 1],
         [1, 0, 0, 0, 1, 2, 0, 2],
         [0, 1, 0, 2, 0, 1, 1, 1],
         [0, 2, 0, 1, 1, 0, 0, 0],
         [2, 0, 1, 1, 1, 0, 0, 2],
         [1, 2, 1, 0, 0, 0, 0, 1]],

        [[2, 0, 0, 2, 2, 2, 1, 2],
         [2, 2, 1, 1, 0, 1, 1, 0],
         [2, 2, 2, 0, 0, 1, 2, 2],
         [2, 2, 2, 0, 1, 1, 1, 1],
         [2, 0, 0, 0, 1, 0, 2, 2],
         [2, 1, 0, 1, 1, 0, 0, 2],
         [1, 2, 1, 1, 0, 0, 1, 2],
         [2, 0, 2, 1, 2, 1, 0, 1]]],


       [[[2, 1, 1, 1, 0, 0, 1, 1],
         [0, 1, 2, 2, 2, 0, 0, 0],
         [1, 2, 0, 2, 0, 0, 2, 2],
         [1, 0, 1, 2, 1, 0, 1, 2],
         [0, 0, 0, 2, 1, 2, 1, 1],
         [0, 1, 2, 2, 0, 0, 1, 2],
         [0, 0, 2, 0, 1, 0, 2, 2],
         [1, 1, 1, 1, 2, 1, 0, 2]],

        [[1, 0, 2, 0, 2, 0, 0, 1],
         [1, 0, 0, 0, 0, 2, 1, 2],
         [1, 0, 1, 0, 2, 0, 2, 1],
         [0, 1, 0, 0, 0, 0, 2, 1],
         [0, 0, 1, 1, 2, 2, 1, 1],
         [0, 2, 1, 1, 0, 0, 0, 2],
         [1, 1, 1, 2, 1, 2, 2, 0],
         [0, 2, 1, 0, 1, 2, 0, 0]],

        [[2, 1, 1, 0, 1, 0, 1, 1],
         [0, 1, 2, 1, 1, 0, 2, 1],
         [1, 1, 0, 0, 2, 1, 1, 1],
         [2, 1, 1, 0, 2, 1, 1, 1],
         [1, 0, 1, 0, 1, 2, 1, 1],
         [0, 2, 2, 0, 0, 0, 0, 0],
         [1, 0, 1, 2, 2, 1, 0, 1],
         [1, 0, 1, 2, 1, 2, 2, 1]],

        [[0, 1, 2, 0, 2, 2, 2, 0],
         [0, 2, 0, 1, 1, 0, 2, 1],
         [0, 2, 2, 2, 0, 1, 2, 2],
         [1, 1, 2, 0, 0, 2, 2, 0],
         [2, 1, 1, 2, 0, 0, 1, 2],
         [1, 2, 1, 1, 2, 2, 2, 0],
         [0, 2, 2, 2, 0, 2, 0, 1],
         [2, 2, 2, 1, 1, 0, 1, 1]]]], dtype=uint8)


*/


//                  W  H  C  N
//reg [`DWIDTH-1:0] a[8][8][4][2] =
//                  N  C  H  W
reg [`DWIDTH-1:0] a[2][4][8][8] =
'{     '{'{'{8'd1, 8'd1, 8'd1, 8'd1, 8'd1, 8'd1, 8'd2, 8'd0},
         '{8'd0, 8'd1, 8'd1, 8'd1, 8'd1, 8'd2, 8'd2, 8'd1},
         '{8'd0, 8'd0, 8'd0, 8'd2, 8'd2, 8'd0, 8'd0, 8'd2},
         '{8'd1, 8'd0, 8'd0, 8'd2, 8'd2, 8'd2, 8'd0, 8'd1},
         '{8'd2, 8'd2, 8'd2, 8'd2, 8'd0, 8'd2, 8'd1, 8'd1},
         '{8'd2, 8'd1, 8'd1, 8'd2, 8'd2, 8'd1, 8'd0, 8'd0},
         '{8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd1, 8'd2, 8'd2},
         '{8'd0, 8'd2, 8'd0, 8'd2, 8'd1, 8'd0, 8'd2, 8'd1}},

        '{'{8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0, 8'd1, 8'd0},
         '{8'd1, 8'd2, 8'd1, 8'd0, 8'd1, 8'd2, 8'd1, 8'd0},
         '{8'd1, 8'd1, 8'd2, 8'd0, 8'd0, 8'd1, 8'd0, 8'd0},
         '{8'd2, 8'd2, 8'd2, 8'd0, 8'd2, 8'd2, 8'd1, 8'd2},
         '{8'd1, 8'd2, 8'd0, 8'd2, 8'd1, 8'd2, 8'd1, 8'd0},
         '{8'd2, 8'd2, 8'd0, 8'd0, 8'd0, 8'd0, 8'd1, 8'd2},
         '{8'd1, 8'd0, 8'd2, 8'd1, 8'd1, 8'd0, 8'd1, 8'd0},
         '{8'd1, 8'd1, 8'd0, 8'd2, 8'd0, 8'd2, 8'd1, 8'd2}},

        '{'{8'd0, 8'd1, 8'd2, 8'd2, 8'd1, 8'd0, 8'd2, 8'd0},
         '{8'd2, 8'd0, 8'd1, 8'd1, 8'd2, 8'd0, 8'd0, 8'd2},
         '{8'd1, 8'd1, 8'd1, 8'd0, 8'd1, 8'd0, 8'd1, 8'd1},
         '{8'd1, 8'd0, 8'd0, 8'd0, 8'd1, 8'd2, 8'd0, 8'd2},
         '{8'd0, 8'd1, 8'd0, 8'd2, 8'd0, 8'd1, 8'd1, 8'd1},
         '{8'd0, 8'd2, 8'd0, 8'd1, 8'd1, 8'd0, 8'd0, 8'd0},
         '{8'd2, 8'd0, 8'd1, 8'd1, 8'd1, 8'd0, 8'd0, 8'd2},
         '{8'd1, 8'd2, 8'd1, 8'd0, 8'd0, 8'd0, 8'd0, 8'd1}},

        '{'{8'd2, 8'd0, 8'd0, 8'd2, 8'd2, 8'd2, 8'd1, 8'd2},
         '{8'd2, 8'd2, 8'd1, 8'd1, 8'd0, 8'd1, 8'd1, 8'd0},
         '{8'd2, 8'd2, 8'd2, 8'd0, 8'd0, 8'd1, 8'd2, 8'd2},
         '{8'd2, 8'd2, 8'd2, 8'd0, 8'd1, 8'd1, 8'd1, 8'd1},
         '{8'd2, 8'd0, 8'd0, 8'd0, 8'd1, 8'd0, 8'd2, 8'd2},
         '{8'd2, 8'd1, 8'd0, 8'd1, 8'd1, 8'd0, 8'd0, 8'd2},
         '{8'd1, 8'd2, 8'd1, 8'd1, 8'd0, 8'd0, 8'd1, 8'd2},
         '{8'd2, 8'd0, 8'd2, 8'd1, 8'd2, 8'd1, 8'd0, 8'd1}}},


       '{'{'{8'd2, 8'd1, 8'd1, 8'd1, 8'd0, 8'd0, 8'd1, 8'd1},
         '{8'd0, 8'd1, 8'd2, 8'd2, 8'd2, 8'd0, 8'd0, 8'd0},
         '{8'd1, 8'd2, 8'd0, 8'd2, 8'd0, 8'd0, 8'd2, 8'd2},
         '{8'd1, 8'd0, 8'd1, 8'd2, 8'd1, 8'd0, 8'd1, 8'd2},
         '{8'd0, 8'd0, 8'd0, 8'd2, 8'd1, 8'd2, 8'd1, 8'd1},
         '{8'd0, 8'd1, 8'd2, 8'd2, 8'd0, 8'd0, 8'd1, 8'd2},
         '{8'd0, 8'd0, 8'd2, 8'd0, 8'd1, 8'd0, 8'd2, 8'd2},
         '{8'd1, 8'd1, 8'd1, 8'd1, 8'd2, 8'd1, 8'd0, 8'd2}},

        '{'{8'd1, 8'd0, 8'd2, 8'd0, 8'd2, 8'd0, 8'd0, 8'd1},
         '{8'd1, 8'd0, 8'd0, 8'd0, 8'd0, 8'd2, 8'd1, 8'd2},
         '{8'd1, 8'd0, 8'd1, 8'd0, 8'd2, 8'd0, 8'd2, 8'd1},
         '{8'd0, 8'd1, 8'd0, 8'd0, 8'd0, 8'd0, 8'd2, 8'd1},
         '{8'd0, 8'd0, 8'd1, 8'd1, 8'd2, 8'd2, 8'd1, 8'd1},
         '{8'd0, 8'd2, 8'd1, 8'd1, 8'd0, 8'd0, 8'd0, 8'd2},
         '{8'd1, 8'd1, 8'd1, 8'd2, 8'd1, 8'd2, 8'd2, 8'd0},
         '{8'd0, 8'd2, 8'd1, 8'd0, 8'd1, 8'd2, 8'd0, 8'd0}},

        '{'{8'd2, 8'd1, 8'd1, 8'd0, 8'd1, 8'd0, 8'd1, 8'd1},
         '{8'd0, 8'd1, 8'd2, 8'd1, 8'd1, 8'd0, 8'd2, 8'd1},
         '{8'd1, 8'd1, 8'd0, 8'd0, 8'd2, 8'd1, 8'd1, 8'd1},
         '{8'd2, 8'd1, 8'd1, 8'd0, 8'd2, 8'd1, 8'd1, 8'd1},
         '{8'd1, 8'd0, 8'd1, 8'd0, 8'd1, 8'd2, 8'd1, 8'd1},
         '{8'd0, 8'd2, 8'd2, 8'd0, 8'd0, 8'd0, 8'd0, 8'd0},
         '{8'd1, 8'd0, 8'd1, 8'd2, 8'd2, 8'd1, 8'd0, 8'd1},
         '{8'd1, 8'd0, 8'd1, 8'd2, 8'd1, 8'd2, 8'd2, 8'd1}},

        '{'{8'd0, 8'd1, 8'd2, 8'd0, 8'd2, 8'd2, 8'd2, 8'd0},
         '{8'd0, 8'd2, 8'd0, 8'd1, 8'd1, 8'd0, 8'd2, 8'd1},
         '{8'd0, 8'd2, 8'd2, 8'd2, 8'd0, 8'd1, 8'd2, 8'd2},
         '{8'd1, 8'd1, 8'd2, 8'd0, 8'd0, 8'd2, 8'd2, 8'd0},
         '{8'd2, 8'd1, 8'd1, 8'd2, 8'd0, 8'd0, 8'd1, 8'd2},
         '{8'd1, 8'd2, 8'd1, 8'd1, 8'd2, 8'd2, 8'd2, 8'd0},
         '{8'd0, 8'd2, 8'd2, 8'd2, 8'd0, 8'd2, 8'd0, 8'd1},
         '{8'd2, 8'd2, 8'd2, 8'd1, 8'd1, 8'd0, 8'd1, 8'd1}}}};



////////////////////////////////////////////
// 4D weights matrix
////////////////////////////////////////////
/*
>>> b = np.random.randint(low=0, high=3,size=(4,4,2,2), dtype=np.uint8)
>>> b
array([[[[1, 0],
         [2, 0]],

        [[2, 0],
         [1, 1]],

        [[0, 2],
         [1, 2]],

        [[0, 0],
         [0, 0]]],


       [[[2, 1],
         [2, 2]],

        [[2, 0],
         [1, 0]],

        [[0, 2],
         [0, 0]],

        [[2, 0],
         [2, 1]]],


       [[[0, 2],
         [1, 0]],

        [[0, 2],
         [0, 1]],

        [[2, 2],
         [2, 2]],

        [[1, 1],
         [0, 1]]],


       [[[2, 0],
         [1, 2]],

        [[1, 1],
         [2, 2]],

        [[2, 2],
         [2, 0]],

        [[0, 0],
         [2, 2]]]], dtype=uint8)

*/
//                  W  H  C  K
//reg [`DWIDTH-1:0] b[2][2][4][4] =
//                  K  C  H  W
reg [`DWIDTH-1:0] b[4][4][2][2] =
'{     '{'{'{8'd1, 8'd0},
         '{8'd2, 8'd0}},

        '{'{8'd2, 8'd0},
         '{8'd1, 8'd1}},

        '{'{8'd0, 8'd2},
         '{8'd1, 8'd2}},

        '{'{8'd0, 8'd0},
         '{8'd0, 8'd0}}},


       '{'{'{8'd2, 8'd1},
         '{8'd2, 8'd2}},

        '{'{8'd2, 8'd0},
         '{8'd1, 8'd0}},

        '{'{8'd0, 8'd2},
         '{8'd0, 8'd0}},

        '{'{8'd2, 8'd0},
         '{8'd2, 8'd1}}},


       '{'{'{8'd0, 8'd2},
         '{8'd1, 8'd0}},

        '{'{8'd0, 8'd2},
         '{8'd0, 8'd1}},

        '{'{8'd2, 8'd2},
         '{8'd2, 8'd2}},

        '{'{8'd1, 8'd1},
         '{8'd0, 8'd1}}},


       '{'{'{8'd2, 8'd0},
         '{8'd1, 8'd2}},

        '{'{8'd1, 8'd1},
         '{8'd2, 8'd2}},

        '{'{8'd2, 8'd2},
         '{8'd2, 8'd0}},

        '{'{8'd0, 8'd0},
         '{8'd2, 8'd2}}}};

////////////////////////////////////////////
//Task to initialize BRAMs
////////////////////////////////////////////
task initialize_brams();
begin
    for (int n=0; n<batch_size; n++) begin
        for (int c=0; c<inp_channels; c++) begin
            for (int h=0; h<inp_height; h++) begin
                for (int w=0; w<inp_width; w++) begin
                    u_top.matrix_A.ram[
                        a_start_addr +
                        n * inp_channels * inp_height * inp_width +
                        c * inp_height * inp_width +
                        h * inp_width +
                        w
                    ] = a[n][c][h][w];
                end
            end    
        end
    end

    for (int n=0; n<out_channels; n++) begin
        for (int c=0; c<inp_channels; c++) begin
            for (int h=0; h<filter_height; h++) begin
                for (int w=0; w<filter_width; w++) begin
                    u_top.matrix_B.ram[
                        b_start_addr +
                        n * inp_channels * filter_height * filter_width +
                        c * filter_height * filter_width +
                        h * filter_width +
                        w
                    ] = b[n][c][h][w];
                end
            end    
        end
    end

end
endtask

////////////////////////////////////////////
//Task to compare outputs with expected values
////////////////////////////////////////////
task compare_outputs();
begin

end
endtask

////////////////////////////////////////////
//The actual test
////////////////////////////////////////////
task convolution_test();
begin
  
end
endtask

endmodule
